module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127;
  wire n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023;
  assign n136 = x125 | x128;
  assign n137 = x126 | x128;
  assign n138 = (x125 & ~n136) | (x125 & n137) | (~n136 & n137);
  assign n139 = x129 & n138;
  assign n140 = x0 | x128;
  assign n141 = (x127 & ~x128) | (x127 & n140) | (~x128 & n140);
  assign n142 = n140 & n141;
  assign n143 = x129 & n142;
  assign n144 = (n139 & n142) | (n139 & ~n143) | (n142 & ~n143);
  assign n145 = (x130 & ~x131) | (x130 & n144) | (~x131 & n144);
  assign n146 = x121 & x128;
  assign n147 = (x122 & ~x128) | (x122 & n146) | (~x128 & n146);
  assign n148 = n146 | n147;
  assign n149 = x129 & n148;
  assign n150 = x123 & x128;
  assign n151 = (x124 & ~x128) | (x124 & n150) | (~x128 & n150);
  assign n152 = n150 | n151;
  assign n153 = x129 & n152;
  assign n154 = (n149 & n152) | (n149 & ~n153) | (n152 & ~n153);
  assign n155 = (x130 & x131) | (x130 & ~n154) | (x131 & ~n154);
  assign n156 = n145 & ~n155;
  assign n157 = ~x118 & x128;
  assign n158 = ~x117 & x128;
  assign n159 = (x118 & n157) | (x118 & ~n158) | (n157 & ~n158);
  assign n160 = x129 & n159;
  assign n161 = x119 & x128;
  assign n162 = (x120 & ~x128) | (x120 & n161) | (~x128 & n161);
  assign n163 = n161 | n162;
  assign n164 = x129 & n163;
  assign n165 = (n160 & n163) | (n160 & ~n164) | (n163 & ~n164);
  assign n166 = (x130 & x131) | (x130 & n165) | (x131 & n165);
  assign n167 = ~x114 & x128;
  assign n168 = ~x113 & x128;
  assign n169 = (x114 & n167) | (x114 & ~n168) | (n167 & ~n168);
  assign n170 = x129 & n169;
  assign n171 = x115 | x128;
  assign n172 = x116 | x128;
  assign n173 = (x115 & ~n171) | (x115 & n172) | (~n171 & n172);
  assign n174 = x129 & n173;
  assign n175 = (n170 & n173) | (n170 & ~n174) | (n173 & ~n174);
  assign n176 = (~x130 & x131) | (~x130 & n175) | (x131 & n175);
  assign n177 = n166 & n176;
  assign n178 = n156 | n177;
  assign n179 = (x132 & ~x133) | (x132 & n178) | (~x133 & n178);
  assign n180 = x109 & x128;
  assign n181 = (x110 & ~x128) | (x110 & n180) | (~x128 & n180);
  assign n182 = n180 | n181;
  assign n183 = x129 & n182;
  assign n184 = x111 & x128;
  assign n185 = (x112 & ~x128) | (x112 & n184) | (~x128 & n184);
  assign n186 = n184 | n185;
  assign n187 = x129 & n186;
  assign n188 = (n183 & n186) | (n183 & ~n187) | (n186 & ~n187);
  assign n189 = (x130 & ~x131) | (x130 & n188) | (~x131 & n188);
  assign n190 = x105 & x128;
  assign n191 = (x106 & ~x128) | (x106 & n190) | (~x128 & n190);
  assign n192 = n190 | n191;
  assign n193 = x129 & n192;
  assign n194 = x107 & x128;
  assign n195 = (x108 & ~x128) | (x108 & n194) | (~x128 & n194);
  assign n196 = n194 | n195;
  assign n197 = x129 & n196;
  assign n198 = (n193 & n196) | (n193 & ~n197) | (n196 & ~n197);
  assign n199 = (x130 & x131) | (x130 & ~n198) | (x131 & ~n198);
  assign n200 = n189 & ~n199;
  assign n201 = x101 & x128;
  assign n202 = (x102 & ~x128) | (x102 & n201) | (~x128 & n201);
  assign n203 = n201 | n202;
  assign n204 = x129 & n203;
  assign n205 = x103 & x128;
  assign n206 = (x104 & ~x128) | (x104 & n205) | (~x128 & n205);
  assign n207 = n205 | n206;
  assign n208 = x129 & n207;
  assign n209 = (n204 & n207) | (n204 & ~n208) | (n207 & ~n208);
  assign n210 = (x130 & x131) | (x130 & n209) | (x131 & n209);
  assign n211 = x97 & x128;
  assign n212 = (x98 & ~x128) | (x98 & n211) | (~x128 & n211);
  assign n213 = n211 | n212;
  assign n214 = x129 & n213;
  assign n215 = x99 & x128;
  assign n216 = (x100 & ~x128) | (x100 & n215) | (~x128 & n215);
  assign n217 = n215 | n216;
  assign n218 = x129 & n217;
  assign n219 = (n214 & n217) | (n214 & ~n218) | (n217 & ~n218);
  assign n220 = (~x130 & x131) | (~x130 & n219) | (x131 & n219);
  assign n221 = n210 & n220;
  assign n222 = n200 | n221;
  assign n223 = (x132 & x133) | (x132 & ~n222) | (x133 & ~n222);
  assign n224 = n179 & ~n223;
  assign n225 = x93 & x128;
  assign n226 = (x94 & ~x128) | (x94 & n225) | (~x128 & n225);
  assign n227 = n225 | n226;
  assign n228 = x129 & n227;
  assign n229 = x95 & x128;
  assign n230 = (x96 & ~x128) | (x96 & n229) | (~x128 & n229);
  assign n231 = n229 | n230;
  assign n232 = x129 & n231;
  assign n233 = (n228 & n231) | (n228 & ~n232) | (n231 & ~n232);
  assign n234 = (x130 & ~x131) | (x130 & n233) | (~x131 & n233);
  assign n235 = x89 & x128;
  assign n236 = (x90 & ~x128) | (x90 & n235) | (~x128 & n235);
  assign n237 = n235 | n236;
  assign n238 = x129 & n237;
  assign n239 = x91 & x128;
  assign n240 = (x92 & ~x128) | (x92 & n239) | (~x128 & n239);
  assign n241 = n239 | n240;
  assign n242 = x129 & n241;
  assign n243 = (n238 & n241) | (n238 & ~n242) | (n241 & ~n242);
  assign n244 = (x130 & x131) | (x130 & ~n243) | (x131 & ~n243);
  assign n245 = n234 & ~n244;
  assign n246 = x85 & x128;
  assign n247 = (x86 & ~x128) | (x86 & n246) | (~x128 & n246);
  assign n248 = n246 | n247;
  assign n249 = x129 & n248;
  assign n250 = x87 & x128;
  assign n251 = (x88 & ~x128) | (x88 & n250) | (~x128 & n250);
  assign n252 = n250 | n251;
  assign n253 = x129 & n252;
  assign n254 = (n249 & n252) | (n249 & ~n253) | (n252 & ~n253);
  assign n255 = (x130 & x131) | (x130 & n254) | (x131 & n254);
  assign n256 = x81 & x128;
  assign n257 = (x82 & ~x128) | (x82 & n256) | (~x128 & n256);
  assign n258 = n256 | n257;
  assign n259 = x129 & n258;
  assign n260 = x83 & x128;
  assign n261 = (x84 & ~x128) | (x84 & n260) | (~x128 & n260);
  assign n262 = n260 | n261;
  assign n263 = x129 & n262;
  assign n264 = (n259 & n262) | (n259 & ~n263) | (n262 & ~n263);
  assign n265 = (~x130 & x131) | (~x130 & n264) | (x131 & n264);
  assign n266 = n255 & n265;
  assign n267 = n245 | n266;
  assign n268 = (x132 & x133) | (x132 & n267) | (x133 & n267);
  assign n269 = x77 & x128;
  assign n270 = (x78 & ~x128) | (x78 & n269) | (~x128 & n269);
  assign n271 = n269 | n270;
  assign n272 = x129 & n271;
  assign n273 = x79 & x128;
  assign n274 = (x80 & ~x128) | (x80 & n273) | (~x128 & n273);
  assign n275 = n273 | n274;
  assign n276 = x129 & n275;
  assign n277 = (n272 & n275) | (n272 & ~n276) | (n275 & ~n276);
  assign n278 = (x130 & ~x131) | (x130 & n277) | (~x131 & n277);
  assign n279 = x73 & x128;
  assign n280 = (x74 & ~x128) | (x74 & n279) | (~x128 & n279);
  assign n281 = n279 | n280;
  assign n282 = x129 & n281;
  assign n283 = x75 & x128;
  assign n284 = (x76 & ~x128) | (x76 & n283) | (~x128 & n283);
  assign n285 = n283 | n284;
  assign n286 = x129 & n285;
  assign n287 = (n282 & n285) | (n282 & ~n286) | (n285 & ~n286);
  assign n288 = (x130 & x131) | (x130 & ~n287) | (x131 & ~n287);
  assign n289 = n278 & ~n288;
  assign n290 = x69 & x128;
  assign n291 = (x70 & ~x128) | (x70 & n290) | (~x128 & n290);
  assign n292 = n290 | n291;
  assign n293 = x129 & n292;
  assign n294 = x71 & x128;
  assign n295 = (x72 & ~x128) | (x72 & n294) | (~x128 & n294);
  assign n296 = n294 | n295;
  assign n297 = x129 & n296;
  assign n298 = (n293 & n296) | (n293 & ~n297) | (n296 & ~n297);
  assign n299 = (x130 & x131) | (x130 & n298) | (x131 & n298);
  assign n300 = x65 & x128;
  assign n301 = (x66 & ~x128) | (x66 & n300) | (~x128 & n300);
  assign n302 = n300 | n301;
  assign n303 = x129 & n302;
  assign n304 = x67 & x128;
  assign n305 = (x68 & ~x128) | (x68 & n304) | (~x128 & n304);
  assign n306 = n304 | n305;
  assign n307 = x129 & n306;
  assign n308 = (n303 & n306) | (n303 & ~n307) | (n306 & ~n307);
  assign n309 = (~x130 & x131) | (~x130 & n308) | (x131 & n308);
  assign n310 = n299 & n309;
  assign n311 = n289 | n310;
  assign n312 = (~x132 & x133) | (~x132 & n311) | (x133 & n311);
  assign n313 = n268 & n312;
  assign n314 = n224 | n313;
  assign n315 = x45 & x128;
  assign n316 = (x46 & ~x128) | (x46 & n315) | (~x128 & n315);
  assign n317 = n315 | n316;
  assign n318 = x129 & n317;
  assign n319 = ~x48 & x128;
  assign n320 = ~x47 & x128;
  assign n321 = (x48 & n319) | (x48 & ~n320) | (n319 & ~n320);
  assign n322 = x129 & n321;
  assign n323 = (n318 & n321) | (n318 & ~n322) | (n321 & ~n322);
  assign n324 = (x130 & ~x131) | (x130 & n323) | (~x131 & n323);
  assign n325 = x41 & x128;
  assign n326 = (x42 & ~x128) | (x42 & n325) | (~x128 & n325);
  assign n327 = n325 | n326;
  assign n328 = x129 & n327;
  assign n329 = x43 | x128;
  assign n330 = x44 | x128;
  assign n331 = (x43 & ~n329) | (x43 & n330) | (~n329 & n330);
  assign n332 = x129 & n331;
  assign n333 = (n328 & n331) | (n328 & ~n332) | (n331 & ~n332);
  assign n334 = (x130 & x131) | (x130 & ~n333) | (x131 & ~n333);
  assign n335 = n324 & ~n334;
  assign n336 = x128 & ~x129;
  assign n337 = ~x39 & x128;
  assign n338 = (x38 & x128) | (x38 & ~x129) | (x128 & ~x129);
  assign n339 = x38 & ~n338;
  assign n340 = (n336 & ~n337) | (n336 & n339) | (~n337 & n339);
  assign n341 = x128 | x129;
  assign n342 = x40 | x128;
  assign n343 = x37 & x129;
  assign n344 = x128 & n343;
  assign n345 = (~n341 & n342) | (~n341 & n344) | (n342 & n344);
  assign n346 = n340 | n345;
  assign n347 = (x130 & x131) | (x130 & n346) | (x131 & n346);
  assign n348 = x33 & x128;
  assign n349 = (x34 & ~x128) | (x34 & n348) | (~x128 & n348);
  assign n350 = n348 | n349;
  assign n351 = x129 & n350;
  assign n352 = x35 & x128;
  assign n353 = (x36 & ~x128) | (x36 & n352) | (~x128 & n352);
  assign n354 = n352 | n353;
  assign n355 = x129 & n354;
  assign n356 = (n351 & n354) | (n351 & ~n355) | (n354 & ~n355);
  assign n357 = (~x130 & x131) | (~x130 & n356) | (x131 & n356);
  assign n358 = n347 & n357;
  assign n359 = n335 | n358;
  assign n360 = (x132 & x133) | (x132 & ~n359) | (x133 & ~n359);
  assign n361 = x61 & x128;
  assign n362 = (x62 & ~x128) | (x62 & n361) | (~x128 & n361);
  assign n363 = n361 | n362;
  assign n364 = x129 & n363;
  assign n365 = x63 & x128;
  assign n366 = (x64 & ~x128) | (x64 & n365) | (~x128 & n365);
  assign n367 = n365 | n366;
  assign n368 = x129 & n367;
  assign n369 = (n364 & n367) | (n364 & ~n368) | (n367 & ~n368);
  assign n370 = (x130 & ~x131) | (x130 & n369) | (~x131 & n369);
  assign n371 = x57 & x128;
  assign n372 = (x58 & ~x128) | (x58 & n371) | (~x128 & n371);
  assign n373 = n371 | n372;
  assign n374 = x129 & n373;
  assign n375 = x59 & x128;
  assign n376 = (x60 & ~x128) | (x60 & n375) | (~x128 & n375);
  assign n377 = n375 | n376;
  assign n378 = x129 & n377;
  assign n379 = (n374 & n377) | (n374 & ~n378) | (n377 & ~n378);
  assign n380 = (x130 & x131) | (x130 & ~n379) | (x131 & ~n379);
  assign n381 = n370 & ~n380;
  assign n382 = x53 & x128;
  assign n383 = (x54 & ~x128) | (x54 & n382) | (~x128 & n382);
  assign n384 = n382 | n383;
  assign n385 = x129 & n384;
  assign n386 = x55 & x128;
  assign n387 = (x56 & ~x128) | (x56 & n386) | (~x128 & n386);
  assign n388 = n386 | n387;
  assign n389 = x129 & n388;
  assign n390 = (n385 & n388) | (n385 & ~n389) | (n388 & ~n389);
  assign n391 = (x130 & x131) | (x130 & n390) | (x131 & n390);
  assign n392 = x49 | x128;
  assign n393 = x50 | x128;
  assign n394 = (x49 & ~n392) | (x49 & n393) | (~n392 & n393);
  assign n395 = x129 & n394;
  assign n396 = x51 & x128;
  assign n397 = (x52 & ~x128) | (x52 & n396) | (~x128 & n396);
  assign n398 = n396 | n397;
  assign n399 = x129 & n398;
  assign n400 = (n395 & n398) | (n395 & ~n399) | (n398 & ~n399);
  assign n401 = (~x130 & x131) | (~x130 & n400) | (x131 & n400);
  assign n402 = n391 & n401;
  assign n403 = n381 | n402;
  assign n404 = (x132 & ~x133) | (x132 & n403) | (~x133 & n403);
  assign n405 = ~n360 & n404;
  assign n406 = x133 | n405;
  assign n407 = x29 & x128;
  assign n408 = (x30 & ~x128) | (x30 & n407) | (~x128 & n407);
  assign n409 = n407 | n408;
  assign n410 = x129 & n409;
  assign n411 = x31 & x128;
  assign n412 = (x32 & ~x128) | (x32 & n411) | (~x128 & n411);
  assign n413 = n411 | n412;
  assign n414 = x129 & n413;
  assign n415 = (n410 & n413) | (n410 & ~n414) | (n413 & ~n414);
  assign n416 = (x130 & ~x131) | (x130 & n415) | (~x131 & n415);
  assign n417 = x25 & x128;
  assign n418 = (x26 & ~x128) | (x26 & n417) | (~x128 & n417);
  assign n419 = n417 | n418;
  assign n420 = x129 & n419;
  assign n421 = x27 & x128;
  assign n422 = (x28 & ~x128) | (x28 & n421) | (~x128 & n421);
  assign n423 = n421 | n422;
  assign n424 = x129 & n423;
  assign n425 = (n420 & n423) | (n420 & ~n424) | (n423 & ~n424);
  assign n426 = (x130 & x131) | (x130 & ~n425) | (x131 & ~n425);
  assign n427 = n416 & ~n426;
  assign n428 = x21 & x128;
  assign n429 = (x22 & ~x128) | (x22 & n428) | (~x128 & n428);
  assign n430 = n428 | n429;
  assign n431 = x129 & n430;
  assign n432 = x23 & x128;
  assign n433 = (x24 & ~x128) | (x24 & n432) | (~x128 & n432);
  assign n434 = n432 | n433;
  assign n435 = x129 & n434;
  assign n436 = (n431 & n434) | (n431 & ~n435) | (n434 & ~n435);
  assign n437 = (x130 & x131) | (x130 & n436) | (x131 & n436);
  assign n438 = x17 & x128;
  assign n439 = (x18 & ~x128) | (x18 & n438) | (~x128 & n438);
  assign n440 = n438 | n439;
  assign n441 = x129 & n440;
  assign n442 = x19 & x128;
  assign n443 = (x20 & ~x128) | (x20 & n442) | (~x128 & n442);
  assign n444 = n442 | n443;
  assign n445 = x129 & n444;
  assign n446 = (n441 & n444) | (n441 & ~n445) | (n444 & ~n445);
  assign n447 = (~x130 & x131) | (~x130 & n446) | (x131 & n446);
  assign n448 = n437 & n447;
  assign n449 = n427 | n448;
  assign n450 = x13 & x128;
  assign n451 = (x14 & ~x128) | (x14 & n450) | (~x128 & n450);
  assign n452 = n450 | n451;
  assign n453 = x129 & n452;
  assign n454 = x15 & x128;
  assign n455 = (x16 & ~x128) | (x16 & n454) | (~x128 & n454);
  assign n456 = n454 | n455;
  assign n457 = x129 & n456;
  assign n458 = (n453 & n456) | (n453 & ~n457) | (n456 & ~n457);
  assign n459 = (x130 & ~x131) | (x130 & n458) | (~x131 & n458);
  assign n460 = x9 & x128;
  assign n461 = (x10 & ~x128) | (x10 & n460) | (~x128 & n460);
  assign n462 = n460 | n461;
  assign n463 = x129 & n462;
  assign n464 = x11 & x128;
  assign n465 = (x12 & ~x128) | (x12 & n464) | (~x128 & n464);
  assign n466 = n464 | n465;
  assign n467 = x129 & n466;
  assign n468 = (n463 & n466) | (n463 & ~n467) | (n466 & ~n467);
  assign n469 = (x130 & x131) | (x130 & ~n468) | (x131 & ~n468);
  assign n470 = n459 & ~n469;
  assign n471 = x5 & x128;
  assign n472 = (x6 & ~x128) | (x6 & n471) | (~x128 & n471);
  assign n473 = n471 | n472;
  assign n474 = x129 & n473;
  assign n475 = x7 & x128;
  assign n476 = (x8 & ~x128) | (x8 & n475) | (~x128 & n475);
  assign n477 = n475 | n476;
  assign n478 = x129 & n477;
  assign n479 = (n474 & n477) | (n474 & ~n478) | (n477 & ~n478);
  assign n480 = (x130 & x131) | (x130 & n479) | (x131 & n479);
  assign n481 = ~x2 & x128;
  assign n482 = ~x1 & x128;
  assign n483 = (x2 & n481) | (x2 & ~n482) | (n481 & ~n482);
  assign n484 = x129 & n483;
  assign n485 = x3 & x128;
  assign n486 = (x4 & ~x128) | (x4 & n485) | (~x128 & n485);
  assign n487 = n485 | n486;
  assign n488 = x129 & n487;
  assign n489 = (n484 & n487) | (n484 & ~n488) | (n487 & ~n488);
  assign n490 = (~x130 & x131) | (~x130 & n489) | (x131 & n489);
  assign n491 = n480 & n490;
  assign n492 = n470 | n491;
  assign n493 = (x132 & ~x133) | (x132 & n492) | (~x133 & n492);
  assign n494 = (~x132 & n449) | (~x132 & n493) | (n449 & n493);
  assign n495 = (n405 & n406) | (n405 & n493) | (n406 & n493);
  assign n496 = (n406 & n494) | (n406 & n495) | (n494 & n495);
  assign n497 = x134 & ~n496;
  assign n498 = x134 & ~n314;
  assign n499 = (n314 & ~n497) | (n314 & n498) | (~n497 & n498);
  assign n500 = x0 & n336;
  assign n501 = (x127 & ~x128) | (x127 & n336) | (~x128 & n336);
  assign n502 = n336 | n501;
  assign n503 = (x129 & n500) | (x129 & n502) | (n500 & n502);
  assign n504 = x1 | x129;
  assign n505 = (x126 & x128) | (x126 & ~n341) | (x128 & ~n341);
  assign n506 = x129 & n505;
  assign n507 = (~n341 & n504) | (~n341 & n506) | (n504 & n506);
  assign n508 = n503 | n507;
  assign n509 = (x130 & ~x131) | (x130 & n508) | (~x131 & n508);
  assign n510 = x124 & n336;
  assign n511 = (x123 & x129) | (x123 & n336) | (x129 & n336);
  assign n512 = n336 | n511;
  assign n513 = (~x128 & n510) | (~x128 & n512) | (n510 & n512);
  assign n514 = (x122 & x129) | (x122 & ~n341) | (x129 & ~n341);
  assign n515 = x128 & n514;
  assign n516 = (n136 & ~n341) | (n136 & n515) | (~n341 & n515);
  assign n517 = n513 | n516;
  assign n518 = (x130 & x131) | (x130 & ~n517) | (x131 & ~n517);
  assign n519 = n509 & ~n518;
  assign n520 = x120 & n336;
  assign n521 = (x119 & x129) | (x119 & n336) | (x129 & n336);
  assign n522 = n336 | n521;
  assign n523 = (~x128 & n520) | (~x128 & n522) | (n520 & n522);
  assign n524 = x121 | x128;
  assign n525 = (x118 & x129) | (x118 & ~n341) | (x129 & ~n341);
  assign n526 = x128 & n525;
  assign n527 = (~n341 & n524) | (~n341 & n526) | (n524 & n526);
  assign n528 = n523 | n527;
  assign n529 = (x130 & x131) | (x130 & n528) | (x131 & n528);
  assign n530 = x114 & x128;
  assign n531 = (x117 & ~x129) | (x117 & n530) | (~x129 & n530);
  assign n532 = n530 | n531;
  assign n533 = n336 & n532;
  assign n534 = x116 & ~x129;
  assign n535 = x115 & ~x128;
  assign n536 = n341 & n535;
  assign n537 = (n341 & n534) | (n341 & n536) | (n534 & n536);
  assign n538 = (n532 & ~n533) | (n532 & n537) | (~n533 & n537);
  assign n539 = (~x130 & x131) | (~x130 & n538) | (x131 & n538);
  assign n540 = n529 & n539;
  assign n541 = n519 | n540;
  assign n542 = (x132 & ~x133) | (x132 & n541) | (~x133 & n541);
  assign n543 = x112 & n336;
  assign n544 = (x111 & x129) | (x111 & n336) | (x129 & n336);
  assign n545 = n336 | n544;
  assign n546 = (~x128 & n543) | (~x128 & n545) | (n543 & n545);
  assign n547 = x113 | x128;
  assign n548 = (x110 & x129) | (x110 & ~n341) | (x129 & ~n341);
  assign n549 = x128 & n548;
  assign n550 = (~n341 & n547) | (~n341 & n549) | (n547 & n549);
  assign n551 = n546 | n550;
  assign n552 = (x130 & ~x131) | (x130 & n551) | (~x131 & n551);
  assign n553 = x108 & n336;
  assign n554 = (x107 & x129) | (x107 & n336) | (x129 & n336);
  assign n555 = n336 | n554;
  assign n556 = (~x128 & n553) | (~x128 & n555) | (n553 & n555);
  assign n557 = x109 | x128;
  assign n558 = (x106 & x129) | (x106 & ~n341) | (x129 & ~n341);
  assign n559 = x128 & n558;
  assign n560 = (~n341 & n557) | (~n341 & n559) | (n557 & n559);
  assign n561 = n556 | n560;
  assign n562 = (x130 & x131) | (x130 & ~n561) | (x131 & ~n561);
  assign n563 = n552 & ~n562;
  assign n564 = x104 & n336;
  assign n565 = (x103 & x129) | (x103 & n336) | (x129 & n336);
  assign n566 = n336 | n565;
  assign n567 = (~x128 & n564) | (~x128 & n566) | (n564 & n566);
  assign n568 = x105 | x128;
  assign n569 = (x102 & x129) | (x102 & ~n341) | (x129 & ~n341);
  assign n570 = x128 & n569;
  assign n571 = (~n341 & n568) | (~n341 & n570) | (n568 & n570);
  assign n572 = n567 | n571;
  assign n573 = (x130 & x131) | (x130 & n572) | (x131 & n572);
  assign n574 = x100 & n336;
  assign n575 = (x99 & x129) | (x99 & n336) | (x129 & n336);
  assign n576 = n336 | n575;
  assign n577 = (~x128 & n574) | (~x128 & n576) | (n574 & n576);
  assign n578 = x101 | x128;
  assign n579 = (x98 & x129) | (x98 & ~n341) | (x129 & ~n341);
  assign n580 = x128 & n579;
  assign n581 = (~n341 & n578) | (~n341 & n580) | (n578 & n580);
  assign n582 = n577 | n581;
  assign n583 = (~x130 & x131) | (~x130 & n582) | (x131 & n582);
  assign n584 = n573 & n583;
  assign n585 = n563 | n584;
  assign n586 = (x132 & x133) | (x132 & ~n585) | (x133 & ~n585);
  assign n587 = n542 & ~n586;
  assign n588 = x96 & n336;
  assign n589 = (x95 & x129) | (x95 & n336) | (x129 & n336);
  assign n590 = n336 | n589;
  assign n591 = (~x128 & n588) | (~x128 & n590) | (n588 & n590);
  assign n592 = x97 | x128;
  assign n593 = (x94 & x129) | (x94 & ~n341) | (x129 & ~n341);
  assign n594 = x128 & n593;
  assign n595 = (~n341 & n592) | (~n341 & n594) | (n592 & n594);
  assign n596 = n591 | n595;
  assign n597 = (x130 & ~x131) | (x130 & n596) | (~x131 & n596);
  assign n598 = x92 & n336;
  assign n599 = (x91 & x129) | (x91 & n336) | (x129 & n336);
  assign n600 = n336 | n599;
  assign n601 = (~x128 & n598) | (~x128 & n600) | (n598 & n600);
  assign n602 = x93 | x128;
  assign n603 = (x90 & x129) | (x90 & ~n341) | (x129 & ~n341);
  assign n604 = x128 & n603;
  assign n605 = (~n341 & n602) | (~n341 & n604) | (n602 & n604);
  assign n606 = n601 | n605;
  assign n607 = (x130 & x131) | (x130 & ~n606) | (x131 & ~n606);
  assign n608 = n597 & ~n607;
  assign n609 = ~x86 & x128;
  assign n610 = x89 & ~x129;
  assign n611 = (x128 & ~n609) | (x128 & n610) | (~n609 & n610);
  assign n612 = ~n336 & n611;
  assign n613 = x88 & n336;
  assign n614 = (x87 & x129) | (x87 & n336) | (x129 & n336);
  assign n615 = n336 | n614;
  assign n616 = (~x128 & n613) | (~x128 & n615) | (n613 & n615);
  assign n617 = n612 | n616;
  assign n618 = (x130 & x131) | (x130 & n617) | (x131 & n617);
  assign n619 = x84 & n336;
  assign n620 = (x83 & x129) | (x83 & n336) | (x129 & n336);
  assign n621 = n336 | n620;
  assign n622 = (~x128 & n619) | (~x128 & n621) | (n619 & n621);
  assign n623 = x85 | x128;
  assign n624 = (x82 & x129) | (x82 & ~n341) | (x129 & ~n341);
  assign n625 = x128 & n624;
  assign n626 = (~n341 & n623) | (~n341 & n625) | (n623 & n625);
  assign n627 = n622 | n626;
  assign n628 = (~x130 & x131) | (~x130 & n627) | (x131 & n627);
  assign n629 = n618 & n628;
  assign n630 = n608 | n629;
  assign n631 = (x132 & x133) | (x132 & n630) | (x133 & n630);
  assign n632 = x80 & n336;
  assign n633 = (x79 & x129) | (x79 & n336) | (x129 & n336);
  assign n634 = n336 | n633;
  assign n635 = (~x128 & n632) | (~x128 & n634) | (n632 & n634);
  assign n636 = x81 | x128;
  assign n637 = (x78 & x129) | (x78 & ~n341) | (x129 & ~n341);
  assign n638 = x128 & n637;
  assign n639 = (~n341 & n636) | (~n341 & n638) | (n636 & n638);
  assign n640 = n635 | n639;
  assign n641 = (x130 & ~x131) | (x130 & n640) | (~x131 & n640);
  assign n642 = x76 & n336;
  assign n643 = (x75 & x129) | (x75 & n336) | (x129 & n336);
  assign n644 = n336 | n643;
  assign n645 = (~x128 & n642) | (~x128 & n644) | (n642 & n644);
  assign n646 = x77 | x128;
  assign n647 = (x74 & x129) | (x74 & ~n341) | (x129 & ~n341);
  assign n648 = x128 & n647;
  assign n649 = (~n341 & n646) | (~n341 & n648) | (n646 & n648);
  assign n650 = n645 | n649;
  assign n651 = (x130 & x131) | (x130 & ~n650) | (x131 & ~n650);
  assign n652 = n641 & ~n651;
  assign n653 = x72 & n336;
  assign n654 = (x71 & x129) | (x71 & n336) | (x129 & n336);
  assign n655 = n336 | n654;
  assign n656 = (~x128 & n653) | (~x128 & n655) | (n653 & n655);
  assign n657 = x73 | x128;
  assign n658 = (x70 & x129) | (x70 & ~n341) | (x129 & ~n341);
  assign n659 = x128 & n658;
  assign n660 = (~n341 & n657) | (~n341 & n659) | (n657 & n659);
  assign n661 = n656 | n660;
  assign n662 = (x130 & x131) | (x130 & n661) | (x131 & n661);
  assign n663 = x68 & n336;
  assign n664 = (x67 & x129) | (x67 & n336) | (x129 & n336);
  assign n665 = n336 | n664;
  assign n666 = (~x128 & n663) | (~x128 & n665) | (n663 & n665);
  assign n667 = x69 | x128;
  assign n668 = (x66 & x129) | (x66 & ~n341) | (x129 & ~n341);
  assign n669 = x128 & n668;
  assign n670 = (~n341 & n667) | (~n341 & n669) | (n667 & n669);
  assign n671 = n666 | n670;
  assign n672 = (~x130 & x131) | (~x130 & n671) | (x131 & n671);
  assign n673 = n662 & n672;
  assign n674 = n652 | n673;
  assign n675 = (~x132 & x133) | (~x132 & n674) | (x133 & n674);
  assign n676 = n631 & n675;
  assign n677 = n587 | n676;
  assign n678 = x132 & ~x133;
  assign n679 = (x47 & x128) | (x47 & ~x129) | (x128 & ~x129);
  assign n680 = x47 & ~n679;
  assign n681 = (~n319 & n336) | (~n319 & n680) | (n336 & n680);
  assign n682 = (~x46 & x128) | (~x46 & x129) | (x128 & x129);
  assign n683 = x46 & n682;
  assign n684 = (~n341 & n392) | (~n341 & n683) | (n392 & n683);
  assign n685 = n681 | n684;
  assign n686 = (x130 & ~x131) | (x130 & n685) | (~x131 & n685);
  assign n687 = x44 & x128;
  assign n688 = (x45 & ~n315) | (x45 & n687) | (~n315 & n687);
  assign n689 = x129 & n688;
  assign n690 = x42 & x128;
  assign n691 = x43 & ~x128;
  assign n692 = (x129 & n690) | (x129 & n691) | (n690 & n691);
  assign n693 = (n688 & ~n689) | (n688 & n692) | (~n689 & n692);
  assign n694 = (x130 & x131) | (x130 & ~n693) | (x131 & ~n693);
  assign n695 = n686 & ~n694;
  assign n696 = (~x40 & x128) | (~x40 & x129) | (x128 & x129);
  assign n697 = (x41 & x128) | (x41 & ~x129) | (x128 & ~x129);
  assign n698 = ~n696 & n697;
  assign n699 = (x39 & x128) | (x39 & x129) | (x128 & x129);
  assign n700 = (x38 & ~x128) | (x38 & x129) | (~x128 & x129);
  assign n701 = n698 | n700;
  assign n702 = (n698 & n699) | (n698 & n701) | (n699 & n701);
  assign n703 = (x130 & x131) | (x130 & n702) | (x131 & n702);
  assign n704 = x36 & n336;
  assign n705 = (x35 & x129) | (x35 & n336) | (x129 & n336);
  assign n706 = n336 | n705;
  assign n707 = (~x128 & n704) | (~x128 & n706) | (n704 & n706);
  assign n708 = x37 | x128;
  assign n709 = (x34 & x129) | (x34 & ~n341) | (x129 & ~n341);
  assign n710 = x128 & n709;
  assign n711 = (~n341 & n708) | (~n341 & n710) | (n708 & n710);
  assign n712 = n707 | n711;
  assign n713 = (~x130 & x131) | (~x130 & n712) | (x131 & n712);
  assign n714 = n703 & n713;
  assign n715 = n695 | n714;
  assign n716 = x133 | n715;
  assign n717 = x32 & n336;
  assign n718 = (x31 & x129) | (x31 & n336) | (x129 & n336);
  assign n719 = n336 | n718;
  assign n720 = (~x128 & n717) | (~x128 & n719) | (n717 & n719);
  assign n721 = x33 | x128;
  assign n722 = (x30 & x129) | (x30 & ~n341) | (x129 & ~n341);
  assign n723 = x128 & n722;
  assign n724 = (~n341 & n721) | (~n341 & n723) | (n721 & n723);
  assign n725 = n720 | n724;
  assign n726 = (x130 & ~x131) | (x130 & n725) | (~x131 & n725);
  assign n727 = x28 & n336;
  assign n728 = (x27 & x129) | (x27 & n336) | (x129 & n336);
  assign n729 = n336 | n728;
  assign n730 = (~x128 & n727) | (~x128 & n729) | (n727 & n729);
  assign n731 = x29 | x128;
  assign n732 = (x26 & x129) | (x26 & ~n341) | (x129 & ~n341);
  assign n733 = x128 & n732;
  assign n734 = (~n341 & n731) | (~n341 & n733) | (n731 & n733);
  assign n735 = n730 | n734;
  assign n736 = (x130 & x131) | (x130 & ~n735) | (x131 & ~n735);
  assign n737 = n726 & ~n736;
  assign n738 = x24 & n336;
  assign n739 = (x23 & x129) | (x23 & n336) | (x129 & n336);
  assign n740 = n336 | n739;
  assign n741 = (~x128 & n738) | (~x128 & n740) | (n738 & n740);
  assign n742 = x25 | x128;
  assign n743 = (x22 & x129) | (x22 & ~n341) | (x129 & ~n341);
  assign n744 = x128 & n743;
  assign n745 = (~n341 & n742) | (~n341 & n744) | (n742 & n744);
  assign n746 = n741 | n745;
  assign n747 = (x130 & x131) | (x130 & n746) | (x131 & n746);
  assign n748 = x20 & n336;
  assign n749 = (x19 & x129) | (x19 & n336) | (x129 & n336);
  assign n750 = n336 | n749;
  assign n751 = (~x128 & n748) | (~x128 & n750) | (n748 & n750);
  assign n752 = x21 | x128;
  assign n753 = (x18 & x129) | (x18 & ~n341) | (x129 & ~n341);
  assign n754 = x128 & n753;
  assign n755 = (~n341 & n752) | (~n341 & n754) | (n752 & n754);
  assign n756 = n751 | n755;
  assign n757 = (~x130 & x131) | (~x130 & n756) | (x131 & n756);
  assign n758 = n747 & n757;
  assign n759 = n737 | n758;
  assign n760 = (x132 & ~x133) | (x132 & n759) | (~x133 & n759);
  assign n761 = n759 & ~n760;
  assign n762 = (n678 & n716) | (n678 & n761) | (n716 & n761);
  assign n763 = x132 | x133;
  assign n764 = x64 & n336;
  assign n765 = (x63 & x129) | (x63 & n336) | (x129 & n336);
  assign n766 = n336 | n765;
  assign n767 = (~x128 & n764) | (~x128 & n766) | (n764 & n766);
  assign n768 = x65 | x128;
  assign n769 = (x62 & x129) | (x62 & ~n341) | (x129 & ~n341);
  assign n770 = x128 & n769;
  assign n771 = (~n341 & n768) | (~n341 & n770) | (n768 & n770);
  assign n772 = n767 | n771;
  assign n773 = (x130 & ~x131) | (x130 & n772) | (~x131 & n772);
  assign n774 = x60 & n336;
  assign n775 = (x59 & x129) | (x59 & n336) | (x129 & n336);
  assign n776 = n336 | n775;
  assign n777 = (~x128 & n774) | (~x128 & n776) | (n774 & n776);
  assign n778 = x61 | x128;
  assign n779 = (x58 & x129) | (x58 & ~n341) | (x129 & ~n341);
  assign n780 = x128 & n779;
  assign n781 = (~n341 & n778) | (~n341 & n780) | (n778 & n780);
  assign n782 = n777 | n781;
  assign n783 = (x130 & x131) | (x130 & ~n782) | (x131 & ~n782);
  assign n784 = n773 & ~n783;
  assign n785 = x56 & n336;
  assign n786 = (x55 & x129) | (x55 & n336) | (x129 & n336);
  assign n787 = n336 | n786;
  assign n788 = (~x128 & n785) | (~x128 & n787) | (n785 & n787);
  assign n789 = x57 | x128;
  assign n790 = (x54 & x129) | (x54 & ~n341) | (x129 & ~n341);
  assign n791 = x128 & n790;
  assign n792 = (~n341 & n789) | (~n341 & n791) | (n789 & n791);
  assign n793 = n788 | n792;
  assign n794 = (x130 & x131) | (x130 & n793) | (x131 & n793);
  assign n795 = x52 & n336;
  assign n796 = (x51 & x129) | (x51 & n336) | (x129 & n336);
  assign n797 = n336 | n796;
  assign n798 = (~x128 & n795) | (~x128 & n797) | (n795 & n797);
  assign n799 = x53 | x128;
  assign n800 = (x50 & x129) | (x50 & ~n341) | (x129 & ~n341);
  assign n801 = x128 & n800;
  assign n802 = (~n341 & n799) | (~n341 & n801) | (n799 & n801);
  assign n803 = n798 | n802;
  assign n804 = (~x130 & x131) | (~x130 & n803) | (x131 & n803);
  assign n805 = n794 & n804;
  assign n806 = n784 | n805;
  assign n807 = x133 | n806;
  assign n808 = x16 & n336;
  assign n809 = (x15 & x129) | (x15 & n336) | (x129 & n336);
  assign n810 = n336 | n809;
  assign n811 = (~x128 & n808) | (~x128 & n810) | (n808 & n810);
  assign n812 = x17 | x128;
  assign n813 = (x14 & x129) | (x14 & ~n341) | (x129 & ~n341);
  assign n814 = x128 & n813;
  assign n815 = (~n341 & n812) | (~n341 & n814) | (n812 & n814);
  assign n816 = n811 | n815;
  assign n817 = (x130 & ~x131) | (x130 & n816) | (~x131 & n816);
  assign n818 = x12 & n336;
  assign n819 = (x11 & x129) | (x11 & n336) | (x129 & n336);
  assign n820 = n336 | n819;
  assign n821 = (~x128 & n818) | (~x128 & n820) | (n818 & n820);
  assign n822 = x13 | x128;
  assign n823 = (x10 & x129) | (x10 & ~n341) | (x129 & ~n341);
  assign n824 = x128 & n823;
  assign n825 = (~n341 & n822) | (~n341 & n824) | (n822 & n824);
  assign n826 = n821 | n825;
  assign n827 = (x130 & x131) | (x130 & ~n826) | (x131 & ~n826);
  assign n828 = n817 & ~n827;
  assign n829 = x8 & n336;
  assign n830 = (x7 & x129) | (x7 & n336) | (x129 & n336);
  assign n831 = n336 | n830;
  assign n832 = (~x128 & n829) | (~x128 & n831) | (n829 & n831);
  assign n833 = x9 | x128;
  assign n834 = (x6 & x129) | (x6 & ~n341) | (x129 & ~n341);
  assign n835 = x128 & n834;
  assign n836 = (~n341 & n833) | (~n341 & n835) | (n833 & n835);
  assign n837 = n832 | n836;
  assign n838 = (x130 & x131) | (x130 & n837) | (x131 & n837);
  assign n839 = x4 & n336;
  assign n840 = (x3 & x129) | (x3 & n336) | (x129 & n336);
  assign n841 = n336 | n840;
  assign n842 = (~x128 & n839) | (~x128 & n841) | (n839 & n841);
  assign n843 = x5 | x128;
  assign n844 = (x2 & x129) | (x2 & ~n341) | (x129 & ~n341);
  assign n845 = x128 & n844;
  assign n846 = (~n341 & n843) | (~n341 & n845) | (n843 & n845);
  assign n847 = n842 | n846;
  assign n848 = (~x130 & x131) | (~x130 & n847) | (x131 & n847);
  assign n849 = n838 & n848;
  assign n850 = n828 | n849;
  assign n851 = (x132 & x133) | (x132 & ~n850) | (x133 & ~n850);
  assign n852 = n850 & n851;
  assign n853 = (~n763 & n807) | (~n763 & n852) | (n807 & n852);
  assign n854 = n762 | n853;
  assign n855 = x134 & ~n854;
  assign n856 = x134 & ~n677;
  assign n857 = (n677 & ~n855) | (n677 & n856) | (~n855 & n856);
  assign n858 = (n143 & n483) | (n143 & ~n484) | (n483 & ~n484);
  assign n859 = (x130 & ~x131) | (x130 & n858) | (~x131 & n858);
  assign n860 = (n138 & ~n139) | (n138 & n153) | (~n139 & n153);
  assign n861 = (x130 & x131) | (x130 & ~n860) | (x131 & ~n860);
  assign n862 = n859 & ~n861;
  assign n863 = (n148 & ~n149) | (n148 & n164) | (~n149 & n164);
  assign n864 = (x130 & x131) | (x130 & n863) | (x131 & n863);
  assign n865 = (n159 & ~n160) | (n159 & n174) | (~n160 & n174);
  assign n866 = (~x130 & x131) | (~x130 & n865) | (x131 & n865);
  assign n867 = n864 & n866;
  assign n868 = n862 | n867;
  assign n869 = (x132 & ~x133) | (x132 & n868) | (~x133 & n868);
  assign n870 = (n169 & ~n170) | (n169 & n187) | (~n170 & n187);
  assign n871 = (x130 & ~x131) | (x130 & n870) | (~x131 & n870);
  assign n872 = (n182 & ~n183) | (n182 & n197) | (~n183 & n197);
  assign n873 = (x130 & x131) | (x130 & ~n872) | (x131 & ~n872);
  assign n874 = n871 & ~n873;
  assign n875 = (n192 & ~n193) | (n192 & n208) | (~n193 & n208);
  assign n876 = (x130 & x131) | (x130 & n875) | (x131 & n875);
  assign n877 = (n203 & ~n204) | (n203 & n218) | (~n204 & n218);
  assign n878 = (~x130 & x131) | (~x130 & n877) | (x131 & n877);
  assign n879 = n876 & n878;
  assign n880 = n874 | n879;
  assign n881 = (x132 & x133) | (x132 & ~n880) | (x133 & ~n880);
  assign n882 = n869 & ~n881;
  assign n883 = (n213 & ~n214) | (n213 & n232) | (~n214 & n232);
  assign n884 = (x130 & ~x131) | (x130 & n883) | (~x131 & n883);
  assign n885 = (n227 & ~n228) | (n227 & n242) | (~n228 & n242);
  assign n886 = (x130 & x131) | (x130 & ~n885) | (x131 & ~n885);
  assign n887 = n884 & ~n886;
  assign n888 = (n237 & ~n238) | (n237 & n253) | (~n238 & n253);
  assign n889 = (x130 & x131) | (x130 & n888) | (x131 & n888);
  assign n890 = (n248 & ~n249) | (n248 & n263) | (~n249 & n263);
  assign n891 = (~x130 & x131) | (~x130 & n890) | (x131 & n890);
  assign n892 = n889 & n891;
  assign n893 = n887 | n892;
  assign n894 = (x132 & x133) | (x132 & n893) | (x133 & n893);
  assign n895 = (n258 & ~n259) | (n258 & n276) | (~n259 & n276);
  assign n896 = (x130 & ~x131) | (x130 & n895) | (~x131 & n895);
  assign n897 = (n271 & ~n272) | (n271 & n286) | (~n272 & n286);
  assign n898 = (x130 & x131) | (x130 & ~n897) | (x131 & ~n897);
  assign n899 = n896 & ~n898;
  assign n900 = (n281 & ~n282) | (n281 & n297) | (~n282 & n297);
  assign n901 = (x130 & x131) | (x130 & n900) | (x131 & n900);
  assign n902 = (n292 & ~n293) | (n292 & n307) | (~n293 & n307);
  assign n903 = (~x130 & x131) | (~x130 & n902) | (x131 & n902);
  assign n904 = n901 & n903;
  assign n905 = n899 | n904;
  assign n906 = (~x132 & x133) | (~x132 & n905) | (x133 & n905);
  assign n907 = n894 & n906;
  assign n908 = n882 | n907;
  assign n909 = (n322 & n394) | (n322 & ~n395) | (n394 & ~n395);
  assign n910 = (x130 & ~x131) | (x130 & n909) | (~x131 & n909);
  assign n911 = (n317 & ~n318) | (n317 & n332) | (~n318 & n332);
  assign n912 = (x130 & x131) | (x130 & ~n911) | (x131 & ~n911);
  assign n913 = n910 & ~n912;
  assign n914 = x39 & x128;
  assign n915 = x40 & ~x128;
  assign n916 = (x129 & n914) | (x129 & n915) | (n914 & n915);
  assign n917 = (n327 & ~n328) | (n327 & n916) | (~n328 & n916);
  assign n918 = (x130 & x131) | (x130 & n917) | (x131 & n917);
  assign n919 = (~x37 & x128) | (~x37 & x129) | (x128 & x129);
  assign n920 = n338 | n355;
  assign n921 = (n355 & ~n919) | (n355 & n920) | (~n919 & n920);
  assign n922 = (~x130 & x131) | (~x130 & n921) | (x131 & n921);
  assign n923 = n918 & n922;
  assign n924 = n913 | n923;
  assign n925 = x133 | n924;
  assign n926 = (n350 & ~n351) | (n350 & n414) | (~n351 & n414);
  assign n927 = (x130 & ~x131) | (x130 & n926) | (~x131 & n926);
  assign n928 = (n409 & ~n410) | (n409 & n424) | (~n410 & n424);
  assign n929 = (x130 & x131) | (x130 & ~n928) | (x131 & ~n928);
  assign n930 = n927 & ~n929;
  assign n931 = (n419 & ~n420) | (n419 & n435) | (~n420 & n435);
  assign n932 = (x130 & x131) | (x130 & n931) | (x131 & n931);
  assign n933 = (n430 & ~n431) | (n430 & n445) | (~n431 & n445);
  assign n934 = (~x130 & x131) | (~x130 & n933) | (x131 & n933);
  assign n935 = n932 & n934;
  assign n936 = n930 | n935;
  assign n937 = (x132 & ~x133) | (x132 & n936) | (~x133 & n936);
  assign n938 = n936 & ~n937;
  assign n939 = (n678 & n925) | (n678 & n938) | (n925 & n938);
  assign n940 = (n302 & ~n303) | (n302 & n368) | (~n303 & n368);
  assign n941 = (x130 & ~x131) | (x130 & n940) | (~x131 & n940);
  assign n942 = (n363 & ~n364) | (n363 & n378) | (~n364 & n378);
  assign n943 = (x130 & x131) | (x130 & ~n942) | (x131 & ~n942);
  assign n944 = n941 & ~n943;
  assign n945 = (n373 & ~n374) | (n373 & n389) | (~n374 & n389);
  assign n946 = (x130 & x131) | (x130 & n945) | (x131 & n945);
  assign n947 = (n384 & ~n385) | (n384 & n399) | (~n385 & n399);
  assign n948 = (~x130 & x131) | (~x130 & n947) | (x131 & n947);
  assign n949 = n946 & n948;
  assign n950 = n944 | n949;
  assign n951 = x133 | n950;
  assign n952 = (n440 & ~n441) | (n440 & n457) | (~n441 & n457);
  assign n953 = (x130 & ~x131) | (x130 & n952) | (~x131 & n952);
  assign n954 = (n452 & ~n453) | (n452 & n467) | (~n453 & n467);
  assign n955 = (x130 & x131) | (x130 & ~n954) | (x131 & ~n954);
  assign n956 = n953 & ~n955;
  assign n957 = (n462 & ~n463) | (n462 & n478) | (~n463 & n478);
  assign n958 = (x130 & x131) | (x130 & n957) | (x131 & n957);
  assign n959 = (n473 & ~n474) | (n473 & n488) | (~n474 & n488);
  assign n960 = (~x130 & x131) | (~x130 & n959) | (x131 & n959);
  assign n961 = n958 & n960;
  assign n962 = n956 | n961;
  assign n963 = (x132 & x133) | (x132 & ~n962) | (x133 & ~n962);
  assign n964 = n962 & n963;
  assign n965 = (~n763 & n951) | (~n763 & n964) | (n951 & n964);
  assign n966 = n939 | n965;
  assign n967 = x134 & ~n966;
  assign n968 = x134 & ~n908;
  assign n969 = (n908 & ~n967) | (n908 & n968) | (~n967 & n968);
  assign n970 = x82 & n336;
  assign n971 = (x81 & x129) | (x81 & n336) | (x129 & n336);
  assign n972 = n336 | n971;
  assign n973 = (~x128 & n970) | (~x128 & n972) | (n970 & n972);
  assign n974 = x83 | x128;
  assign n975 = (x80 & x129) | (x80 & ~n341) | (x129 & ~n341);
  assign n976 = x128 & n975;
  assign n977 = (~n341 & n974) | (~n341 & n976) | (n974 & n976);
  assign n978 = n973 | n977;
  assign n979 = (x130 & ~x131) | (x130 & n978) | (~x131 & n978);
  assign n980 = x78 & n336;
  assign n981 = (x77 & x129) | (x77 & n336) | (x129 & n336);
  assign n982 = n336 | n981;
  assign n983 = (~x128 & n980) | (~x128 & n982) | (n980 & n982);
  assign n984 = x79 | x128;
  assign n985 = (x76 & x129) | (x76 & ~n341) | (x129 & ~n341);
  assign n986 = x128 & n985;
  assign n987 = (~n341 & n984) | (~n341 & n986) | (n984 & n986);
  assign n988 = n983 | n987;
  assign n989 = (x130 & x131) | (x130 & ~n988) | (x131 & ~n988);
  assign n990 = n979 & ~n989;
  assign n991 = x74 & n336;
  assign n992 = (x73 & x129) | (x73 & n336) | (x129 & n336);
  assign n993 = n336 | n992;
  assign n994 = (~x128 & n991) | (~x128 & n993) | (n991 & n993);
  assign n995 = x75 | x128;
  assign n996 = (x72 & x129) | (x72 & ~n341) | (x129 & ~n341);
  assign n997 = x128 & n996;
  assign n998 = (~n341 & n995) | (~n341 & n997) | (n995 & n997);
  assign n999 = n994 | n998;
  assign n1000 = (x130 & x131) | (x130 & n999) | (x131 & n999);
  assign n1001 = x70 & n336;
  assign n1002 = (x69 & x129) | (x69 & n336) | (x129 & n336);
  assign n1003 = n336 | n1002;
  assign n1004 = (~x128 & n1001) | (~x128 & n1003) | (n1001 & n1003);
  assign n1005 = x71 | x128;
  assign n1006 = (x68 & x129) | (x68 & ~n341) | (x129 & ~n341);
  assign n1007 = x128 & n1006;
  assign n1008 = (~n341 & n1005) | (~n341 & n1007) | (n1005 & n1007);
  assign n1009 = n1004 | n1008;
  assign n1010 = (~x130 & x131) | (~x130 & n1009) | (x131 & n1009);
  assign n1011 = n1000 & n1010;
  assign n1012 = n990 | n1011;
  assign n1013 = (x132 & ~x133) | (x132 & n1012) | (~x133 & n1012);
  assign n1014 = x133 & n1013;
  assign n1015 = x1 & x129;
  assign n1016 = ~x128 & n1015;
  assign n1017 = (n336 & ~n481) | (n336 & n1016) | (~n481 & n1016);
  assign n1018 = x3 | x128;
  assign n1019 = (x0 & x129) | (x0 & ~n341) | (x129 & ~n341);
  assign n1020 = x128 & n1019;
  assign n1021 = (~n341 & n1018) | (~n341 & n1020) | (n1018 & n1020);
  assign n1022 = n1017 | n1021;
  assign n1023 = (x130 & ~x131) | (x130 & n1022) | (~x131 & n1022);
  assign n1024 = x126 & ~x129;
  assign n1025 = (~x128 & n136) | (~x128 & n1024) | (n136 & n1024);
  assign n1026 = n341 & n1025;
  assign n1027 = x127 | x128;
  assign n1028 = (x124 & x129) | (x124 & ~n341) | (x129 & ~n341);
  assign n1029 = x128 & n1028;
  assign n1030 = (~n341 & n1027) | (~n341 & n1029) | (n1027 & n1029);
  assign n1031 = n1026 | n1030;
  assign n1032 = (x130 & x131) | (x130 & ~n1031) | (x131 & ~n1031);
  assign n1033 = n1023 & ~n1032;
  assign n1034 = x122 & n336;
  assign n1035 = (x121 & x129) | (x121 & n336) | (x129 & n336);
  assign n1036 = n336 | n1035;
  assign n1037 = (~x128 & n1034) | (~x128 & n1036) | (n1034 & n1036);
  assign n1038 = x123 | x128;
  assign n1039 = (x120 & x129) | (x120 & ~n341) | (x129 & ~n341);
  assign n1040 = x128 & n1039;
  assign n1041 = (~n341 & n1038) | (~n341 & n1040) | (n1038 & n1040);
  assign n1042 = n1037 | n1041;
  assign n1043 = (x130 & x131) | (x130 & n1042) | (x131 & n1042);
  assign n1044 = x117 & x129;
  assign n1045 = ~x128 & n1044;
  assign n1046 = (~n157 & n336) | (~n157 & n1045) | (n336 & n1045);
  assign n1047 = x119 | x128;
  assign n1048 = (x116 & x129) | (x116 & ~n341) | (x129 & ~n341);
  assign n1049 = x128 & n1048;
  assign n1050 = (~n341 & n1047) | (~n341 & n1049) | (n1047 & n1049);
  assign n1051 = n1046 | n1050;
  assign n1052 = (~x130 & x131) | (~x130 & n1051) | (x131 & n1051);
  assign n1053 = n1043 & n1052;
  assign n1054 = n1033 | n1053;
  assign n1055 = x133 | n1054;
  assign n1056 = (~n763 & n1014) | (~n763 & n1055) | (n1014 & n1055);
  assign n1057 = x106 & n336;
  assign n1058 = (x105 & x129) | (x105 & n336) | (x129 & n336);
  assign n1059 = n336 | n1058;
  assign n1060 = (~x128 & n1057) | (~x128 & n1059) | (n1057 & n1059);
  assign n1061 = x107 | x128;
  assign n1062 = (x104 & x129) | (x104 & ~n341) | (x129 & ~n341);
  assign n1063 = x128 & n1062;
  assign n1064 = (~n341 & n1061) | (~n341 & n1063) | (n1061 & n1063);
  assign n1065 = n1060 | n1064;
  assign n1066 = (x130 & x131) | (x130 & n1065) | (x131 & n1065);
  assign n1067 = x112 & x128;
  assign n1068 = x129 & n1067;
  assign n1069 = (n171 & ~n341) | (n171 & n1068) | (~n341 & n1068);
  assign n1070 = x113 & x129;
  assign n1071 = ~x128 & n1070;
  assign n1072 = (~n167 & n336) | (~n167 & n1071) | (n336 & n1071);
  assign n1073 = n1069 | n1072;
  assign n1074 = (x130 & ~x131) | (x130 & n1073) | (~x131 & n1073);
  assign n1075 = x110 & n336;
  assign n1076 = (x109 & x129) | (x109 & n336) | (x129 & n336);
  assign n1077 = n336 | n1076;
  assign n1078 = (~x128 & n1075) | (~x128 & n1077) | (n1075 & n1077);
  assign n1079 = x111 | x128;
  assign n1080 = (x108 & x129) | (x108 & ~n341) | (x129 & ~n341);
  assign n1081 = x128 & n1080;
  assign n1082 = (~n341 & n1079) | (~n341 & n1081) | (n1079 & n1081);
  assign n1083 = n1078 | n1082;
  assign n1084 = (x130 & x131) | (x130 & ~n1083) | (x131 & ~n1083);
  assign n1085 = n1074 & ~n1084;
  assign n1086 = x102 & n336;
  assign n1087 = (x101 & x129) | (x101 & n336) | (x129 & n336);
  assign n1088 = n336 | n1087;
  assign n1089 = (~x128 & n1086) | (~x128 & n1088) | (n1086 & n1088);
  assign n1090 = x103 | x128;
  assign n1091 = (x100 & x129) | (x100 & ~n341) | (x129 & ~n341);
  assign n1092 = x128 & n1091;
  assign n1093 = (~n341 & n1090) | (~n341 & n1092) | (n1090 & n1092);
  assign n1094 = n1089 | n1093;
  assign n1095 = (~x130 & x131) | (~x130 & n1094) | (x131 & n1094);
  assign n1096 = n1066 & ~n1095;
  assign n1097 = (n1066 & n1085) | (n1066 & ~n1096) | (n1085 & ~n1096);
  assign n1098 = x133 | n1097;
  assign n1099 = x90 & n336;
  assign n1100 = (x89 & x129) | (x89 & n336) | (x129 & n336);
  assign n1101 = n336 | n1100;
  assign n1102 = (~x128 & n1099) | (~x128 & n1101) | (n1099 & n1101);
  assign n1103 = x91 | x128;
  assign n1104 = (x88 & x129) | (x88 & ~n341) | (x129 & ~n341);
  assign n1105 = x128 & n1104;
  assign n1106 = (~n341 & n1103) | (~n341 & n1105) | (n1103 & n1105);
  assign n1107 = n1102 | n1106;
  assign n1108 = (x130 & x131) | (x130 & n1107) | (x131 & n1107);
  assign n1109 = x98 & n336;
  assign n1110 = (x97 & x129) | (x97 & n336) | (x129 & n336);
  assign n1111 = n336 | n1110;
  assign n1112 = (~x128 & n1109) | (~x128 & n1111) | (n1109 & n1111);
  assign n1113 = x99 | x128;
  assign n1114 = (x96 & x129) | (x96 & ~n341) | (x129 & ~n341);
  assign n1115 = x128 & n1114;
  assign n1116 = (~n341 & n1113) | (~n341 & n1115) | (n1113 & n1115);
  assign n1117 = n1112 | n1116;
  assign n1118 = (x130 & ~x131) | (x130 & n1117) | (~x131 & n1117);
  assign n1119 = x94 & n336;
  assign n1120 = (x93 & x129) | (x93 & n336) | (x129 & n336);
  assign n1121 = n336 | n1120;
  assign n1122 = (~x128 & n1119) | (~x128 & n1121) | (n1119 & n1121);
  assign n1123 = x95 | x128;
  assign n1124 = (x92 & x129) | (x92 & ~n341) | (x129 & ~n341);
  assign n1125 = x128 & n1124;
  assign n1126 = (~n341 & n1123) | (~n341 & n1125) | (n1123 & n1125);
  assign n1127 = n1122 | n1126;
  assign n1128 = (x130 & x131) | (x130 & ~n1127) | (x131 & ~n1127);
  assign n1129 = n1118 & ~n1128;
  assign n1130 = x85 & x129;
  assign n1131 = ~x128 & n1130;
  assign n1132 = (n336 & ~n609) | (n336 & n1131) | (~n609 & n1131);
  assign n1133 = x87 | x128;
  assign n1134 = (x84 & x129) | (x84 & ~n341) | (x129 & ~n341);
  assign n1135 = x128 & n1134;
  assign n1136 = (~n341 & n1133) | (~n341 & n1135) | (n1133 & n1135);
  assign n1137 = n1132 | n1136;
  assign n1138 = (~x130 & x131) | (~x130 & n1137) | (x131 & n1137);
  assign n1139 = n1108 & ~n1138;
  assign n1140 = (n1108 & n1129) | (n1108 & ~n1139) | (n1129 & ~n1139);
  assign n1141 = (x133 & n678) | (x133 & n1140) | (n678 & n1140);
  assign n1142 = ~x132 & n1141;
  assign n1143 = (n678 & n1098) | (n678 & n1142) | (n1098 & n1142);
  assign n1144 = n1056 | n1143;
  assign n1145 = x34 & n336;
  assign n1146 = (x33 & x129) | (x33 & n336) | (x129 & n336);
  assign n1147 = n336 | n1146;
  assign n1148 = (~x128 & n1145) | (~x128 & n1147) | (n1145 & n1147);
  assign n1149 = x35 | x128;
  assign n1150 = (x32 & x129) | (x32 & ~n341) | (x129 & ~n341);
  assign n1151 = x128 & n1150;
  assign n1152 = (~n341 & n1149) | (~n341 & n1151) | (n1149 & n1151);
  assign n1153 = n1148 | n1152;
  assign n1154 = (x130 & ~x131) | (x130 & n1153) | (~x131 & n1153);
  assign n1155 = x30 & n336;
  assign n1156 = (x29 & x129) | (x29 & n336) | (x129 & n336);
  assign n1157 = n336 | n1156;
  assign n1158 = (~x128 & n1155) | (~x128 & n1157) | (n1155 & n1157);
  assign n1159 = x31 | x128;
  assign n1160 = (x28 & x129) | (x28 & ~n341) | (x129 & ~n341);
  assign n1161 = x128 & n1160;
  assign n1162 = (~n341 & n1159) | (~n341 & n1161) | (n1159 & n1161);
  assign n1163 = n1158 | n1162;
  assign n1164 = (x130 & x131) | (x130 & ~n1163) | (x131 & ~n1163);
  assign n1165 = n1154 & ~n1164;
  assign n1166 = x26 & n336;
  assign n1167 = (x25 & x129) | (x25 & n336) | (x129 & n336);
  assign n1168 = n336 | n1167;
  assign n1169 = (~x128 & n1166) | (~x128 & n1168) | (n1166 & n1168);
  assign n1170 = x27 | x128;
  assign n1171 = (x24 & x129) | (x24 & ~n341) | (x129 & ~n341);
  assign n1172 = x128 & n1171;
  assign n1173 = (~n341 & n1170) | (~n341 & n1172) | (n1170 & n1172);
  assign n1174 = n1169 | n1173;
  assign n1175 = (x130 & x131) | (x130 & n1174) | (x131 & n1174);
  assign n1176 = x22 & n336;
  assign n1177 = (x21 & x129) | (x21 & n336) | (x129 & n336);
  assign n1178 = n336 | n1177;
  assign n1179 = (~x128 & n1176) | (~x128 & n1178) | (n1176 & n1178);
  assign n1180 = x23 | x128;
  assign n1181 = (x20 & x129) | (x20 & ~n341) | (x129 & ~n341);
  assign n1182 = x128 & n1181;
  assign n1183 = (~n341 & n1180) | (~n341 & n1182) | (n1180 & n1182);
  assign n1184 = n1179 | n1183;
  assign n1185 = (~x130 & x131) | (~x130 & n1184) | (x131 & n1184);
  assign n1186 = n1175 & n1185;
  assign n1187 = n1165 | n1186;
  assign n1188 = (x132 & x133) | (x132 & n1187) | (x133 & n1187);
  assign n1189 = x18 & n336;
  assign n1190 = (x17 & x129) | (x17 & n336) | (x129 & n336);
  assign n1191 = n336 | n1190;
  assign n1192 = (~x128 & n1189) | (~x128 & n1191) | (n1189 & n1191);
  assign n1193 = x19 | x128;
  assign n1194 = (x16 & x129) | (x16 & ~n341) | (x129 & ~n341);
  assign n1195 = x128 & n1194;
  assign n1196 = (~n341 & n1193) | (~n341 & n1195) | (n1193 & n1195);
  assign n1197 = n1192 | n1196;
  assign n1198 = (x130 & ~x131) | (x130 & n1197) | (~x131 & n1197);
  assign n1199 = x14 & n336;
  assign n1200 = (x13 & x129) | (x13 & n336) | (x129 & n336);
  assign n1201 = n336 | n1200;
  assign n1202 = (~x128 & n1199) | (~x128 & n1201) | (n1199 & n1201);
  assign n1203 = x15 | x128;
  assign n1204 = (x12 & x129) | (x12 & ~n341) | (x129 & ~n341);
  assign n1205 = x128 & n1204;
  assign n1206 = (~n341 & n1203) | (~n341 & n1205) | (n1203 & n1205);
  assign n1207 = n1202 | n1206;
  assign n1208 = (x130 & x131) | (x130 & ~n1207) | (x131 & ~n1207);
  assign n1209 = n1198 & ~n1208;
  assign n1210 = x10 & n336;
  assign n1211 = (x9 & x129) | (x9 & n336) | (x129 & n336);
  assign n1212 = n336 | n1211;
  assign n1213 = (~x128 & n1210) | (~x128 & n1212) | (n1210 & n1212);
  assign n1214 = x11 | x128;
  assign n1215 = (x8 & x129) | (x8 & ~n341) | (x129 & ~n341);
  assign n1216 = x128 & n1215;
  assign n1217 = (~n341 & n1214) | (~n341 & n1216) | (n1214 & n1216);
  assign n1218 = n1213 | n1217;
  assign n1219 = (x130 & x131) | (x130 & n1218) | (x131 & n1218);
  assign n1220 = x6 & n336;
  assign n1221 = (x5 & x129) | (x5 & n336) | (x129 & n336);
  assign n1222 = n336 | n1221;
  assign n1223 = (~x128 & n1220) | (~x128 & n1222) | (n1220 & n1222);
  assign n1224 = x7 | x128;
  assign n1225 = (x4 & x129) | (x4 & ~n341) | (x129 & ~n341);
  assign n1226 = x128 & n1225;
  assign n1227 = (~n341 & n1224) | (~n341 & n1226) | (n1224 & n1226);
  assign n1228 = n1223 | n1227;
  assign n1229 = (~x130 & x131) | (~x130 & n1228) | (x131 & n1228);
  assign n1230 = n1219 & n1229;
  assign n1231 = n1209 | n1230;
  assign n1232 = (~x132 & x133) | (~x132 & n1231) | (x133 & n1231);
  assign n1233 = n1188 & n1232;
  assign n1234 = x50 & n336;
  assign n1235 = (x49 & x129) | (x49 & n336) | (x129 & n336);
  assign n1236 = n336 | n1235;
  assign n1237 = (~x128 & n1234) | (~x128 & n1236) | (n1234 & n1236);
  assign n1238 = x51 | x128;
  assign n1239 = (x48 & x129) | (x48 & ~n341) | (x129 & ~n341);
  assign n1240 = x128 & n1239;
  assign n1241 = (~n341 & n1238) | (~n341 & n1240) | (n1238 & n1240);
  assign n1242 = n1237 | n1241;
  assign n1243 = (x130 & ~x131) | (x130 & n1242) | (~x131 & n1242);
  assign n1244 = (n679 & ~n682) | (n679 & n689) | (~n682 & n689);
  assign n1245 = n689 | n1244;
  assign n1246 = (x130 & x131) | (x130 & ~n1245) | (x131 & ~n1245);
  assign n1247 = n1243 & ~n1246;
  assign n1248 = x40 & n696;
  assign n1249 = (n329 & ~n341) | (n329 & n1248) | (~n341 & n1248);
  assign n1250 = ~x42 & x128;
  assign n1251 = x41 & ~n697;
  assign n1252 = (n336 & ~n1250) | (n336 & n1251) | (~n1250 & n1251);
  assign n1253 = n1249 | n1252;
  assign n1254 = (x130 & x131) | (x130 & n1253) | (x131 & n1253);
  assign n1255 = x39 | x128;
  assign n1256 = (x36 & x129) | (x36 & ~n341) | (x129 & ~n341);
  assign n1257 = x128 & n1256;
  assign n1258 = (~n341 & n1255) | (~n341 & n1257) | (n1255 & n1257);
  assign n1259 = x38 & n336;
  assign n1260 = n336 | n343;
  assign n1261 = (~x128 & n1259) | (~x128 & n1260) | (n1259 & n1260);
  assign n1262 = n1258 | n1261;
  assign n1263 = (~x130 & x131) | (~x130 & n1262) | (x131 & n1262);
  assign n1264 = n1254 & n1263;
  assign n1265 = n1247 | n1264;
  assign n1266 = x132 & n1265;
  assign n1267 = x66 & n336;
  assign n1268 = (x65 & x129) | (x65 & n336) | (x129 & n336);
  assign n1269 = n336 | n1268;
  assign n1270 = (~x128 & n1267) | (~x128 & n1269) | (n1267 & n1269);
  assign n1271 = x67 | x128;
  assign n1272 = (x64 & x129) | (x64 & ~n341) | (x129 & ~n341);
  assign n1273 = x128 & n1272;
  assign n1274 = (~n341 & n1271) | (~n341 & n1273) | (n1271 & n1273);
  assign n1275 = n1270 | n1274;
  assign n1276 = x62 & n336;
  assign n1277 = (x61 & x129) | (x61 & n336) | (x129 & n336);
  assign n1278 = n336 | n1277;
  assign n1279 = (~x128 & n1276) | (~x128 & n1278) | (n1276 & n1278);
  assign n1280 = x63 | x128;
  assign n1281 = (x60 & x129) | (x60 & ~n341) | (x129 & ~n341);
  assign n1282 = x128 & n1281;
  assign n1283 = (~n341 & n1280) | (~n341 & n1282) | (n1280 & n1282);
  assign n1284 = n1279 | n1283;
  assign n1285 = (x130 & x131) | (x130 & n1284) | (x131 & n1284);
  assign n1286 = (~x130 & n1275) | (~x130 & n1285) | (n1275 & n1285);
  assign n1287 = x58 & n336;
  assign n1288 = (x57 & x129) | (x57 & n336) | (x129 & n336);
  assign n1289 = n336 | n1288;
  assign n1290 = (~x128 & n1287) | (~x128 & n1289) | (n1287 & n1289);
  assign n1291 = x59 | x128;
  assign n1292 = (x56 & x129) | (x56 & ~n341) | (x129 & ~n341);
  assign n1293 = x128 & n1292;
  assign n1294 = (~n341 & n1291) | (~n341 & n1293) | (n1291 & n1293);
  assign n1295 = n1290 | n1294;
  assign n1296 = (x130 & x131) | (x130 & n1295) | (x131 & n1295);
  assign n1297 = x54 & n336;
  assign n1298 = (x53 & x129) | (x53 & n336) | (x129 & n336);
  assign n1299 = n336 | n1298;
  assign n1300 = (~x128 & n1297) | (~x128 & n1299) | (n1297 & n1299);
  assign n1301 = x55 | x128;
  assign n1302 = (x52 & x129) | (x52 & ~n341) | (x129 & ~n341);
  assign n1303 = x128 & n1302;
  assign n1304 = (~n341 & n1301) | (~n341 & n1303) | (n1301 & n1303);
  assign n1305 = n1300 | n1304;
  assign n1306 = (~x130 & x131) | (~x130 & n1305) | (x131 & n1305);
  assign n1307 = n1296 & n1306;
  assign n1308 = x131 & ~n1307;
  assign n1309 = (n1285 & n1307) | (n1285 & ~n1308) | (n1307 & ~n1308);
  assign n1310 = (n1286 & ~n1308) | (n1286 & n1309) | (~n1308 & n1309);
  assign n1311 = ~x132 & n1310;
  assign n1312 = (~x133 & n1266) | (~x133 & n1311) | (n1266 & n1311);
  assign n1313 = n1233 | n1312;
  assign n1314 = x134 & ~n1313;
  assign n1315 = x134 & ~n1144;
  assign n1316 = (n1144 & ~n1314) | (n1144 & n1315) | (~n1314 & n1315);
  assign n1317 = (~x130 & x131) | (~x130 & n346) | (x131 & n346);
  assign n1318 = x130 & n323;
  assign n1319 = ~x130 & n400;
  assign n1320 = (~x131 & n1318) | (~x131 & n1319) | (n1318 & n1319);
  assign n1321 = (x130 & x131) | (x130 & n333) | (x131 & n333);
  assign n1322 = n1320 | n1321;
  assign n1323 = (n1317 & n1320) | (n1317 & n1322) | (n1320 & n1322);
  assign n1324 = (x132 & x133) | (x132 & ~n1323) | (x133 & ~n1323);
  assign n1325 = (x130 & ~x131) | (x130 & n308) | (~x131 & n308);
  assign n1326 = (x130 & x131) | (x130 & ~n369) | (x131 & ~n369);
  assign n1327 = n1325 & n1326;
  assign n1328 = (x130 & x131) | (x130 & n379) | (x131 & n379);
  assign n1329 = (~x130 & x131) | (~x130 & n390) | (x131 & n390);
  assign n1330 = n1328 & n1329;
  assign n1331 = (n1325 & ~n1327) | (n1325 & n1330) | (~n1327 & n1330);
  assign n1332 = (x132 & ~x133) | (x132 & n1331) | (~x133 & n1331);
  assign n1333 = ~n1324 & n1332;
  assign n1334 = (x130 & ~x131) | (x130 & n446) | (~x131 & n446);
  assign n1335 = (x130 & x131) | (x130 & ~n458) | (x131 & ~n458);
  assign n1336 = n1334 & n1335;
  assign n1337 = (x130 & x131) | (x130 & n468) | (x131 & n468);
  assign n1338 = (~x130 & x131) | (~x130 & n479) | (x131 & n479);
  assign n1339 = n1337 & n1338;
  assign n1340 = (n1334 & ~n1336) | (n1334 & n1339) | (~n1336 & n1339);
  assign n1341 = (~x132 & x133) | (~x132 & n1340) | (x133 & n1340);
  assign n1342 = (x130 & ~x131) | (x130 & n356) | (~x131 & n356);
  assign n1343 = (x130 & x131) | (x130 & ~n415) | (x131 & ~n415);
  assign n1344 = n1342 & n1343;
  assign n1345 = (x130 & x131) | (x130 & n425) | (x131 & n425);
  assign n1346 = (~x130 & x131) | (~x130 & n436) | (x131 & n436);
  assign n1347 = n1345 & n1346;
  assign n1348 = (n1342 & ~n1344) | (n1342 & n1347) | (~n1344 & n1347);
  assign n1349 = (x132 & x133) | (x132 & n1348) | (x133 & n1348);
  assign n1350 = n1333 | n1349;
  assign n1351 = (n1333 & n1341) | (n1333 & n1350) | (n1341 & n1350);
  assign n1352 = x134 & ~n1351;
  assign n1353 = (x130 & ~x131) | (x130 & n219) | (~x131 & n219);
  assign n1354 = (x130 & x131) | (x130 & ~n233) | (x131 & ~n233);
  assign n1355 = n1353 & n1354;
  assign n1356 = (x130 & x131) | (x130 & n243) | (x131 & n243);
  assign n1357 = (~x130 & x131) | (~x130 & n254) | (x131 & n254);
  assign n1358 = n1356 & n1357;
  assign n1359 = (n1353 & ~n1355) | (n1353 & n1358) | (~n1355 & n1358);
  assign n1360 = (x132 & x133) | (x132 & n1359) | (x133 & n1359);
  assign n1361 = (x130 & ~x131) | (x130 & n264) | (~x131 & n264);
  assign n1362 = (x130 & x131) | (x130 & ~n277) | (x131 & ~n277);
  assign n1363 = n1361 & n1362;
  assign n1364 = (x130 & x131) | (x130 & n287) | (x131 & n287);
  assign n1365 = (~x130 & x131) | (~x130 & n298) | (x131 & n298);
  assign n1366 = n1364 & n1365;
  assign n1367 = (n1361 & ~n1363) | (n1361 & n1366) | (~n1363 & n1366);
  assign n1368 = (~x132 & x133) | (~x132 & n1367) | (x133 & n1367);
  assign n1369 = n1360 & n1368;
  assign n1370 = (x130 & ~x131) | (x130 & n175) | (~x131 & n175);
  assign n1371 = (x130 & x131) | (x130 & ~n188) | (x131 & ~n188);
  assign n1372 = n1370 & ~n1371;
  assign n1373 = (x130 & x131) | (x130 & n198) | (x131 & n198);
  assign n1374 = (~x130 & x131) | (~x130 & n209) | (x131 & n209);
  assign n1375 = n1373 & n1374;
  assign n1376 = n1372 | n1375;
  assign n1377 = (x132 & x133) | (x132 & ~n1376) | (x133 & ~n1376);
  assign n1378 = (~x130 & x131) | (~x130 & n165) | (x131 & n165);
  assign n1379 = x130 & n144;
  assign n1380 = ~x130 & n489;
  assign n1381 = (~x131 & n1379) | (~x131 & n1380) | (n1379 & n1380);
  assign n1382 = (x130 & x131) | (x130 & n154) | (x131 & n154);
  assign n1383 = n1381 | n1382;
  assign n1384 = (n1378 & n1381) | (n1378 & n1383) | (n1381 & n1383);
  assign n1385 = (x132 & ~x133) | (x132 & n1384) | (~x133 & n1384);
  assign n1386 = n1369 | n1385;
  assign n1387 = (n1369 & ~n1377) | (n1369 & n1386) | (~n1377 & n1386);
  assign n1388 = x134 & ~n1387;
  assign n1389 = (~n1352 & n1387) | (~n1352 & n1388) | (n1387 & n1388);
  assign n1390 = (~x130 & x131) | (~x130 & n702) | (x131 & n702);
  assign n1391 = x130 & n685;
  assign n1392 = ~x130 & n803;
  assign n1393 = (~x131 & n1391) | (~x131 & n1392) | (n1391 & n1392);
  assign n1394 = (x130 & x131) | (x130 & n693) | (x131 & n693);
  assign n1395 = n1393 | n1394;
  assign n1396 = (n1390 & n1393) | (n1390 & n1395) | (n1393 & n1395);
  assign n1397 = (x132 & x133) | (x132 & ~n1396) | (x133 & ~n1396);
  assign n1398 = (x130 & ~x131) | (x130 & n671) | (~x131 & n671);
  assign n1399 = (x130 & x131) | (x130 & ~n772) | (x131 & ~n772);
  assign n1400 = n1398 & n1399;
  assign n1401 = (x130 & x131) | (x130 & n782) | (x131 & n782);
  assign n1402 = (~x130 & x131) | (~x130 & n793) | (x131 & n793);
  assign n1403 = n1401 & n1402;
  assign n1404 = (n1398 & ~n1400) | (n1398 & n1403) | (~n1400 & n1403);
  assign n1405 = (x132 & ~x133) | (x132 & n1404) | (~x133 & n1404);
  assign n1406 = ~n1397 & n1405;
  assign n1407 = (x130 & ~x131) | (x130 & n756) | (~x131 & n756);
  assign n1408 = (x130 & x131) | (x130 & ~n816) | (x131 & ~n816);
  assign n1409 = n1407 & n1408;
  assign n1410 = (x130 & x131) | (x130 & n826) | (x131 & n826);
  assign n1411 = (~x130 & x131) | (~x130 & n837) | (x131 & n837);
  assign n1412 = n1410 & n1411;
  assign n1413 = (n1407 & ~n1409) | (n1407 & n1412) | (~n1409 & n1412);
  assign n1414 = (~x132 & x133) | (~x132 & n1413) | (x133 & n1413);
  assign n1415 = (x130 & ~x131) | (x130 & n712) | (~x131 & n712);
  assign n1416 = (x130 & x131) | (x130 & ~n725) | (x131 & ~n725);
  assign n1417 = n1415 & n1416;
  assign n1418 = (x130 & x131) | (x130 & n735) | (x131 & n735);
  assign n1419 = (~x130 & x131) | (~x130 & n746) | (x131 & n746);
  assign n1420 = n1418 & n1419;
  assign n1421 = (n1415 & ~n1417) | (n1415 & n1420) | (~n1417 & n1420);
  assign n1422 = (x132 & x133) | (x132 & n1421) | (x133 & n1421);
  assign n1423 = n1406 | n1422;
  assign n1424 = (n1406 & n1414) | (n1406 & n1423) | (n1414 & n1423);
  assign n1425 = x134 & ~n1424;
  assign n1426 = (x130 & ~x131) | (x130 & n582) | (~x131 & n582);
  assign n1427 = (x130 & x131) | (x130 & ~n596) | (x131 & ~n596);
  assign n1428 = n1426 & n1427;
  assign n1429 = (x130 & x131) | (x130 & n606) | (x131 & n606);
  assign n1430 = (~x130 & x131) | (~x130 & n617) | (x131 & n617);
  assign n1431 = n1429 & n1430;
  assign n1432 = (n1426 & ~n1428) | (n1426 & n1431) | (~n1428 & n1431);
  assign n1433 = (x132 & x133) | (x132 & n1432) | (x133 & n1432);
  assign n1434 = (x130 & ~x131) | (x130 & n627) | (~x131 & n627);
  assign n1435 = (x130 & x131) | (x130 & ~n640) | (x131 & ~n640);
  assign n1436 = n1434 & n1435;
  assign n1437 = (x130 & x131) | (x130 & n650) | (x131 & n650);
  assign n1438 = (~x130 & x131) | (~x130 & n661) | (x131 & n661);
  assign n1439 = n1437 & n1438;
  assign n1440 = (n1434 & ~n1436) | (n1434 & n1439) | (~n1436 & n1439);
  assign n1441 = (~x132 & x133) | (~x132 & n1440) | (x133 & n1440);
  assign n1442 = n1433 & n1441;
  assign n1443 = (x130 & ~x131) | (x130 & n538) | (~x131 & n538);
  assign n1444 = (x130 & x131) | (x130 & ~n551) | (x131 & ~n551);
  assign n1445 = n1443 & ~n1444;
  assign n1446 = (x130 & x131) | (x130 & n561) | (x131 & n561);
  assign n1447 = (~x130 & x131) | (~x130 & n572) | (x131 & n572);
  assign n1448 = n1446 & n1447;
  assign n1449 = n1445 | n1448;
  assign n1450 = (x132 & x133) | (x132 & ~n1449) | (x133 & ~n1449);
  assign n1451 = (~x130 & x131) | (~x130 & n528) | (x131 & n528);
  assign n1452 = x130 & n508;
  assign n1453 = ~x130 & n847;
  assign n1454 = (~x131 & n1452) | (~x131 & n1453) | (n1452 & n1453);
  assign n1455 = (x130 & x131) | (x130 & n517) | (x131 & n517);
  assign n1456 = n1454 | n1455;
  assign n1457 = (n1451 & n1454) | (n1451 & n1456) | (n1454 & n1456);
  assign n1458 = (x132 & ~x133) | (x132 & n1457) | (~x133 & n1457);
  assign n1459 = n1442 | n1458;
  assign n1460 = (n1442 & ~n1450) | (n1442 & n1459) | (~n1450 & n1459);
  assign n1461 = x134 & ~n1460;
  assign n1462 = (~n1425 & n1460) | (~n1425 & n1461) | (n1460 & n1461);
  assign n1463 = (~x130 & x131) | (~x130 & n917) | (x131 & n917);
  assign n1464 = x130 & n909;
  assign n1465 = ~x130 & n947;
  assign n1466 = (~x131 & n1464) | (~x131 & n1465) | (n1464 & n1465);
  assign n1467 = (x130 & x131) | (x130 & n911) | (x131 & n911);
  assign n1468 = n1466 | n1467;
  assign n1469 = (n1463 & n1466) | (n1463 & n1468) | (n1466 & n1468);
  assign n1470 = (x132 & x133) | (x132 & ~n1469) | (x133 & ~n1469);
  assign n1471 = (x130 & ~x131) | (x130 & n902) | (~x131 & n902);
  assign n1472 = (x130 & x131) | (x130 & ~n940) | (x131 & ~n940);
  assign n1473 = n1471 & n1472;
  assign n1474 = (x130 & x131) | (x130 & n942) | (x131 & n942);
  assign n1475 = (~x130 & x131) | (~x130 & n945) | (x131 & n945);
  assign n1476 = n1474 & n1475;
  assign n1477 = (n1471 & ~n1473) | (n1471 & n1476) | (~n1473 & n1476);
  assign n1478 = (x132 & ~x133) | (x132 & n1477) | (~x133 & n1477);
  assign n1479 = ~n1470 & n1478;
  assign n1480 = (x130 & ~x131) | (x130 & n933) | (~x131 & n933);
  assign n1481 = (x130 & x131) | (x130 & ~n952) | (x131 & ~n952);
  assign n1482 = n1480 & n1481;
  assign n1483 = (x130 & x131) | (x130 & n954) | (x131 & n954);
  assign n1484 = (~x130 & x131) | (~x130 & n957) | (x131 & n957);
  assign n1485 = n1483 & n1484;
  assign n1486 = (n1480 & ~n1482) | (n1480 & n1485) | (~n1482 & n1485);
  assign n1487 = (~x132 & x133) | (~x132 & n1486) | (x133 & n1486);
  assign n1488 = (x130 & x131) | (x130 & ~n926) | (x131 & ~n926);
  assign n1489 = (x130 & ~x131) | (x130 & n921) | (~x131 & n921);
  assign n1490 = n1488 | n1489;
  assign n1491 = (x130 & x131) | (x130 & n928) | (x131 & n928);
  assign n1492 = (~x130 & x131) | (~x130 & n931) | (x131 & n931);
  assign n1493 = n1491 & n1492;
  assign n1494 = (~n1488 & n1490) | (~n1488 & n1493) | (n1490 & n1493);
  assign n1495 = (x132 & x133) | (x132 & n1494) | (x133 & n1494);
  assign n1496 = n1479 | n1495;
  assign n1497 = (n1479 & n1487) | (n1479 & n1496) | (n1487 & n1496);
  assign n1498 = x134 & ~n1497;
  assign n1499 = (x130 & ~x131) | (x130 & n877) | (~x131 & n877);
  assign n1500 = (x130 & x131) | (x130 & ~n883) | (x131 & ~n883);
  assign n1501 = n1499 & n1500;
  assign n1502 = (x130 & x131) | (x130 & n885) | (x131 & n885);
  assign n1503 = (~x130 & x131) | (~x130 & n888) | (x131 & n888);
  assign n1504 = n1502 & n1503;
  assign n1505 = (n1499 & ~n1501) | (n1499 & n1504) | (~n1501 & n1504);
  assign n1506 = (x132 & x133) | (x132 & n1505) | (x133 & n1505);
  assign n1507 = (x130 & ~x131) | (x130 & n890) | (~x131 & n890);
  assign n1508 = (x130 & x131) | (x130 & ~n895) | (x131 & ~n895);
  assign n1509 = n1507 & n1508;
  assign n1510 = (x130 & x131) | (x130 & n897) | (x131 & n897);
  assign n1511 = (~x130 & x131) | (~x130 & n900) | (x131 & n900);
  assign n1512 = n1510 & n1511;
  assign n1513 = (n1507 & ~n1509) | (n1507 & n1512) | (~n1509 & n1512);
  assign n1514 = (~x132 & x133) | (~x132 & n1513) | (x133 & n1513);
  assign n1515 = n1506 & n1514;
  assign n1516 = (x130 & ~x131) | (x130 & n865) | (~x131 & n865);
  assign n1517 = (x130 & x131) | (x130 & ~n870) | (x131 & ~n870);
  assign n1518 = n1516 & ~n1517;
  assign n1519 = (x130 & x131) | (x130 & n872) | (x131 & n872);
  assign n1520 = (~x130 & x131) | (~x130 & n875) | (x131 & n875);
  assign n1521 = n1519 & n1520;
  assign n1522 = n1518 | n1521;
  assign n1523 = (x132 & x133) | (x132 & ~n1522) | (x133 & ~n1522);
  assign n1524 = (~x130 & x131) | (~x130 & n863) | (x131 & n863);
  assign n1525 = x130 & n858;
  assign n1526 = ~x130 & n959;
  assign n1527 = (~x131 & n1525) | (~x131 & n1526) | (n1525 & n1526);
  assign n1528 = (x130 & x131) | (x130 & n860) | (x131 & n860);
  assign n1529 = n1527 | n1528;
  assign n1530 = (n1524 & n1527) | (n1524 & n1529) | (n1527 & n1529);
  assign n1531 = (x132 & ~x133) | (x132 & n1530) | (~x133 & n1530);
  assign n1532 = n1515 | n1531;
  assign n1533 = (n1515 & ~n1523) | (n1515 & n1532) | (~n1523 & n1532);
  assign n1534 = x134 & ~n1533;
  assign n1535 = (~n1498 & n1533) | (~n1498 & n1534) | (n1533 & n1534);
  assign n1536 = (~x130 & x131) | (~x130 & n1174) | (x131 & n1174);
  assign n1537 = x130 & n1153;
  assign n1538 = ~x130 & n1262;
  assign n1539 = (~x131 & n1537) | (~x131 & n1538) | (n1537 & n1538);
  assign n1540 = (x130 & x131) | (x130 & n1163) | (x131 & n1163);
  assign n1541 = n1539 | n1540;
  assign n1542 = (n1536 & n1539) | (n1536 & n1541) | (n1539 & n1541);
  assign n1543 = (x132 & x133) | (x132 & n1542) | (x133 & n1542);
  assign n1544 = (x130 & ~x131) | (x130 & n1184) | (~x131 & n1184);
  assign n1545 = (x130 & x131) | (x130 & ~n1197) | (x131 & ~n1197);
  assign n1546 = n1544 & n1545;
  assign n1547 = (x130 & x131) | (x130 & n1207) | (x131 & n1207);
  assign n1548 = (~x130 & x131) | (~x130 & n1218) | (x131 & n1218);
  assign n1549 = n1547 & n1548;
  assign n1550 = (n1544 & ~n1546) | (n1544 & n1549) | (~n1546 & n1549);
  assign n1551 = (~x132 & x133) | (~x132 & n1550) | (x133 & n1550);
  assign n1552 = n1543 & n1551;
  assign n1553 = (~x130 & x131) | (~x130 & n1295) | (x131 & n1295);
  assign n1554 = n1285 & n1553;
  assign n1555 = (x130 & x131) | (x130 & ~n1275) | (x131 & ~n1275);
  assign n1556 = (x130 & ~x131) | (x130 & n1009) | (~x131 & n1009);
  assign n1557 = n1554 | n1556;
  assign n1558 = (n1554 & ~n1555) | (n1554 & n1557) | (~n1555 & n1557);
  assign n1559 = (x132 & ~x133) | (x132 & n1558) | (~x133 & n1558);
  assign n1560 = ~x130 & n1305;
  assign n1561 = x130 & x131;
  assign n1562 = (x130 & ~x131) | (x130 & n1253) | (~x131 & n1253);
  assign n1563 = x131 & ~n1562;
  assign n1564 = (n1560 & n1561) | (n1560 & ~n1563) | (n1561 & ~n1563);
  assign n1565 = (x130 & ~x131) | (x130 & n1245) | (~x131 & n1245);
  assign n1566 = n1245 & ~n1565;
  assign n1567 = x130 | x131;
  assign n1568 = ~x131 & n1242;
  assign n1569 = (n1566 & n1567) | (n1566 & n1568) | (n1567 & n1568);
  assign n1570 = n1564 | n1569;
  assign n1571 = (x132 & x133) | (x132 & ~n1570) | (x133 & ~n1570);
  assign n1572 = ~n1552 & n1571;
  assign n1573 = (n1552 & n1559) | (n1552 & ~n1572) | (n1559 & ~n1572);
  assign n1574 = x134 & ~n1573;
  assign n1575 = (x130 & ~x131) | (x130 & n1051) | (~x131 & n1051);
  assign n1576 = (x130 & x131) | (x130 & ~n1073) | (x131 & ~n1073);
  assign n1577 = n1575 & n1576;
  assign n1578 = (x130 & x131) | (x130 & n1083) | (x131 & n1083);
  assign n1579 = (~x130 & x131) | (~x130 & n1065) | (x131 & n1065);
  assign n1580 = n1578 & n1579;
  assign n1581 = (n1575 & ~n1577) | (n1575 & n1580) | (~n1577 & n1580);
  assign n1582 = (x132 & x133) | (x132 & ~n1581) | (x133 & ~n1581);
  assign n1583 = (~x130 & x131) | (~x130 & n1042) | (x131 & n1042);
  assign n1584 = x130 & n1022;
  assign n1585 = ~x130 & n1228;
  assign n1586 = (~x131 & n1584) | (~x131 & n1585) | (n1584 & n1585);
  assign n1587 = (x130 & x131) | (x130 & n1031) | (x131 & n1031);
  assign n1588 = n1586 | n1587;
  assign n1589 = (n1583 & n1586) | (n1583 & n1588) | (n1586 & n1588);
  assign n1590 = (x132 & ~x133) | (x132 & n1589) | (~x133 & n1589);
  assign n1591 = ~n1582 & n1590;
  assign n1592 = (~x130 & x131) | (~x130 & n999) | (x131 & n999);
  assign n1593 = x130 & n978;
  assign n1594 = ~x130 & n1137;
  assign n1595 = (~x131 & n1593) | (~x131 & n1594) | (n1593 & n1594);
  assign n1596 = (x130 & x131) | (x130 & n988) | (x131 & n988);
  assign n1597 = n1595 | n1596;
  assign n1598 = (n1592 & n1595) | (n1592 & n1597) | (n1595 & n1597);
  assign n1599 = (~x132 & x133) | (~x132 & n1598) | (x133 & n1598);
  assign n1600 = (x130 & ~x131) | (x130 & n1094) | (~x131 & n1094);
  assign n1601 = (x130 & x131) | (x130 & ~n1117) | (x131 & ~n1117);
  assign n1602 = n1600 & ~n1601;
  assign n1603 = (x130 & x131) | (x130 & n1127) | (x131 & n1127);
  assign n1604 = (~x130 & x131) | (~x130 & n1107) | (x131 & n1107);
  assign n1605 = n1603 & n1604;
  assign n1606 = n1602 | n1605;
  assign n1607 = (x132 & x133) | (x132 & n1606) | (x133 & n1606);
  assign n1608 = n1599 & ~n1607;
  assign n1609 = (n1591 & n1599) | (n1591 & ~n1608) | (n1599 & ~n1608);
  assign n1610 = x134 & ~n1609;
  assign n1611 = (~n1574 & n1609) | (~n1574 & n1610) | (n1609 & n1610);
  assign n1612 = (x130 & x131) | (x130 & n415) | (x131 & n415);
  assign n1613 = (~x130 & x131) | (~x130 & n425) | (x131 & n425);
  assign n1614 = n1612 & n1613;
  assign n1615 = x130 & n356;
  assign n1616 = ~x130 & n346;
  assign n1617 = (~x131 & n1615) | (~x131 & n1616) | (n1615 & n1616);
  assign n1618 = n1614 | n1617;
  assign n1619 = (x132 & x133) | (x132 & n1618) | (x133 & n1618);
  assign n1620 = (x130 & ~x131) | (x130 & n436) | (~x131 & n436);
  assign n1621 = (x130 & x131) | (x130 & ~n446) | (x131 & ~n446);
  assign n1622 = n1620 & n1621;
  assign n1623 = (x130 & x131) | (x130 & n458) | (x131 & n458);
  assign n1624 = (~x130 & x131) | (~x130 & n468) | (x131 & n468);
  assign n1625 = n1623 & n1624;
  assign n1626 = (n1620 & ~n1622) | (n1620 & n1625) | (~n1622 & n1625);
  assign n1627 = (~x132 & x133) | (~x132 & n1626) | (x133 & n1626);
  assign n1628 = n1619 & n1627;
  assign n1629 = (x130 & ~x131) | (x130 & n298) | (~x131 & n298);
  assign n1630 = (x130 & x131) | (x130 & ~n308) | (x131 & ~n308);
  assign n1631 = n1629 & n1630;
  assign n1632 = (x130 & x131) | (x130 & n369) | (x131 & n369);
  assign n1633 = (~x130 & x131) | (~x130 & n379) | (x131 & n379);
  assign n1634 = n1632 & n1633;
  assign n1635 = (n1629 & ~n1631) | (n1629 & n1634) | (~n1631 & n1634);
  assign n1636 = (x132 & ~x133) | (x132 & n1635) | (~x133 & n1635);
  assign n1637 = (x130 & ~x131) | (x130 & n390) | (~x131 & n390);
  assign n1638 = (x130 & x131) | (x130 & ~n400) | (x131 & ~n400);
  assign n1639 = n1637 & n1638;
  assign n1640 = (x130 & x131) | (x130 & n323) | (x131 & n323);
  assign n1641 = (~x130 & x131) | (~x130 & n333) | (x131 & n333);
  assign n1642 = n1640 & n1641;
  assign n1643 = (n1637 & ~n1639) | (n1637 & n1642) | (~n1639 & n1642);
  assign n1644 = (x132 & x133) | (x132 & ~n1643) | (x133 & ~n1643);
  assign n1645 = ~n1628 & n1644;
  assign n1646 = (n1628 & n1636) | (n1628 & ~n1645) | (n1636 & ~n1645);
  assign n1647 = x134 & ~n1646;
  assign n1648 = (x130 & ~x131) | (x130 & n165) | (~x131 & n165);
  assign n1649 = (x130 & x131) | (x130 & ~n175) | (x131 & ~n175);
  assign n1650 = n1648 & n1649;
  assign n1651 = (x130 & x131) | (x130 & n188) | (x131 & n188);
  assign n1652 = (~x130 & x131) | (~x130 & n198) | (x131 & n198);
  assign n1653 = n1651 & n1652;
  assign n1654 = (n1648 & ~n1650) | (n1648 & n1653) | (~n1650 & n1653);
  assign n1655 = (x132 & x133) | (x132 & ~n1654) | (x133 & ~n1654);
  assign n1656 = (x130 & ~x131) | (x130 & n479) | (~x131 & n479);
  assign n1657 = (x130 & x131) | (x130 & ~n489) | (x131 & ~n489);
  assign n1658 = n1656 & n1657;
  assign n1659 = (x130 & x131) | (x130 & n144) | (x131 & n144);
  assign n1660 = (~x130 & x131) | (~x130 & n154) | (x131 & n154);
  assign n1661 = n1659 & n1660;
  assign n1662 = (n1656 & ~n1658) | (n1656 & n1661) | (~n1658 & n1661);
  assign n1663 = (x132 & ~x133) | (x132 & n1662) | (~x133 & n1662);
  assign n1664 = ~n1655 & n1663;
  assign n1665 = (x130 & ~x131) | (x130 & n254) | (~x131 & n254);
  assign n1666 = (x130 & x131) | (x130 & ~n264) | (x131 & ~n264);
  assign n1667 = n1665 & n1666;
  assign n1668 = (x130 & x131) | (x130 & n277) | (x131 & n277);
  assign n1669 = (~x130 & x131) | (~x130 & n287) | (x131 & n287);
  assign n1670 = n1668 & n1669;
  assign n1671 = (n1665 & ~n1667) | (n1665 & n1670) | (~n1667 & n1670);
  assign n1672 = (~x132 & x133) | (~x132 & n1671) | (x133 & n1671);
  assign n1673 = (x130 & ~x131) | (x130 & n209) | (~x131 & n209);
  assign n1674 = (x130 & x131) | (x130 & ~n219) | (x131 & ~n219);
  assign n1675 = n1673 & n1674;
  assign n1676 = (x130 & x131) | (x130 & n233) | (x131 & n233);
  assign n1677 = (~x130 & x131) | (~x130 & n243) | (x131 & n243);
  assign n1678 = n1676 & n1677;
  assign n1679 = (n1673 & ~n1675) | (n1673 & n1678) | (~n1675 & n1678);
  assign n1680 = (x132 & x133) | (x132 & n1679) | (x133 & n1679);
  assign n1681 = n1672 & ~n1680;
  assign n1682 = (n1664 & n1672) | (n1664 & ~n1681) | (n1672 & ~n1681);
  assign n1683 = x134 & ~n1682;
  assign n1684 = (~n1647 & n1682) | (~n1647 & n1683) | (n1682 & n1683);
  assign n1685 = (x130 & x131) | (x130 & n725) | (x131 & n725);
  assign n1686 = (~x130 & x131) | (~x130 & n735) | (x131 & n735);
  assign n1687 = n1685 & n1686;
  assign n1688 = x130 & n712;
  assign n1689 = ~x130 & n702;
  assign n1690 = (~x131 & n1688) | (~x131 & n1689) | (n1688 & n1689);
  assign n1691 = n1687 | n1690;
  assign n1692 = (x132 & x133) | (x132 & n1691) | (x133 & n1691);
  assign n1693 = (x130 & ~x131) | (x130 & n746) | (~x131 & n746);
  assign n1694 = (x130 & x131) | (x130 & ~n756) | (x131 & ~n756);
  assign n1695 = n1693 & n1694;
  assign n1696 = (x130 & x131) | (x130 & n816) | (x131 & n816);
  assign n1697 = (~x130 & x131) | (~x130 & n826) | (x131 & n826);
  assign n1698 = n1696 & n1697;
  assign n1699 = (n1693 & ~n1695) | (n1693 & n1698) | (~n1695 & n1698);
  assign n1700 = (~x132 & x133) | (~x132 & n1699) | (x133 & n1699);
  assign n1701 = n1692 & n1700;
  assign n1702 = (x130 & ~x131) | (x130 & n661) | (~x131 & n661);
  assign n1703 = (x130 & x131) | (x130 & ~n671) | (x131 & ~n671);
  assign n1704 = n1702 & n1703;
  assign n1705 = (x130 & x131) | (x130 & n772) | (x131 & n772);
  assign n1706 = (~x130 & x131) | (~x130 & n782) | (x131 & n782);
  assign n1707 = n1705 & n1706;
  assign n1708 = (n1702 & ~n1704) | (n1702 & n1707) | (~n1704 & n1707);
  assign n1709 = (x132 & ~x133) | (x132 & n1708) | (~x133 & n1708);
  assign n1710 = (x130 & ~x131) | (x130 & n793) | (~x131 & n793);
  assign n1711 = (x130 & x131) | (x130 & ~n803) | (x131 & ~n803);
  assign n1712 = n1710 & n1711;
  assign n1713 = (x130 & x131) | (x130 & n685) | (x131 & n685);
  assign n1714 = (~x130 & x131) | (~x130 & n693) | (x131 & n693);
  assign n1715 = n1713 & n1714;
  assign n1716 = (n1710 & ~n1712) | (n1710 & n1715) | (~n1712 & n1715);
  assign n1717 = (x132 & x133) | (x132 & ~n1716) | (x133 & ~n1716);
  assign n1718 = ~n1701 & n1717;
  assign n1719 = (n1701 & n1709) | (n1701 & ~n1718) | (n1709 & ~n1718);
  assign n1720 = x134 & ~n1719;
  assign n1721 = (x130 & ~x131) | (x130 & n528) | (~x131 & n528);
  assign n1722 = (x130 & x131) | (x130 & ~n538) | (x131 & ~n538);
  assign n1723 = n1721 & n1722;
  assign n1724 = (x130 & x131) | (x130 & n551) | (x131 & n551);
  assign n1725 = (~x130 & x131) | (~x130 & n561) | (x131 & n561);
  assign n1726 = n1724 & n1725;
  assign n1727 = (n1721 & ~n1723) | (n1721 & n1726) | (~n1723 & n1726);
  assign n1728 = (x132 & x133) | (x132 & ~n1727) | (x133 & ~n1727);
  assign n1729 = (x130 & ~x131) | (x130 & n837) | (~x131 & n837);
  assign n1730 = (x130 & x131) | (x130 & ~n847) | (x131 & ~n847);
  assign n1731 = n1729 & n1730;
  assign n1732 = (x130 & x131) | (x130 & n508) | (x131 & n508);
  assign n1733 = (~x130 & x131) | (~x130 & n517) | (x131 & n517);
  assign n1734 = n1732 & n1733;
  assign n1735 = (n1729 & ~n1731) | (n1729 & n1734) | (~n1731 & n1734);
  assign n1736 = (x132 & ~x133) | (x132 & n1735) | (~x133 & n1735);
  assign n1737 = ~n1728 & n1736;
  assign n1738 = (x130 & ~x131) | (x130 & n617) | (~x131 & n617);
  assign n1739 = (x130 & x131) | (x130 & ~n627) | (x131 & ~n627);
  assign n1740 = n1738 & n1739;
  assign n1741 = (x130 & x131) | (x130 & n640) | (x131 & n640);
  assign n1742 = (~x130 & x131) | (~x130 & n650) | (x131 & n650);
  assign n1743 = n1741 & n1742;
  assign n1744 = (n1738 & ~n1740) | (n1738 & n1743) | (~n1740 & n1743);
  assign n1745 = (~x132 & x133) | (~x132 & n1744) | (x133 & n1744);
  assign n1746 = (x130 & ~x131) | (x130 & n572) | (~x131 & n572);
  assign n1747 = (x130 & x131) | (x130 & ~n582) | (x131 & ~n582);
  assign n1748 = n1746 & n1747;
  assign n1749 = (x130 & x131) | (x130 & n596) | (x131 & n596);
  assign n1750 = (~x130 & x131) | (~x130 & n606) | (x131 & n606);
  assign n1751 = n1749 & n1750;
  assign n1752 = (n1746 & ~n1748) | (n1746 & n1751) | (~n1748 & n1751);
  assign n1753 = (x132 & x133) | (x132 & n1752) | (x133 & n1752);
  assign n1754 = n1745 & ~n1753;
  assign n1755 = (n1737 & n1745) | (n1737 & ~n1754) | (n1745 & ~n1754);
  assign n1756 = x134 & ~n1755;
  assign n1757 = (~n1720 & n1755) | (~n1720 & n1756) | (n1755 & n1756);
  assign n1758 = (x130 & ~x131) | (x130 & n957) | (~x131 & n957);
  assign n1759 = (x130 & x131) | (x130 & ~n959) | (x131 & ~n959);
  assign n1760 = n1758 & n1759;
  assign n1761 = (x130 & x131) | (x130 & n858) | (x131 & n858);
  assign n1762 = (~x130 & x131) | (~x130 & n860) | (x131 & n860);
  assign n1763 = n1761 & n1762;
  assign n1764 = (n1758 & ~n1760) | (n1758 & n1763) | (~n1760 & n1763);
  assign n1765 = (x132 & ~x133) | (x132 & n1764) | (~x133 & n1764);
  assign n1766 = (x130 & ~x131) | (x130 & n863) | (~x131 & n863);
  assign n1767 = (x130 & x131) | (x130 & ~n865) | (x131 & ~n865);
  assign n1768 = n1766 & n1767;
  assign n1769 = (x130 & x131) | (x130 & n870) | (x131 & n870);
  assign n1770 = (~x130 & x131) | (~x130 & n872) | (x131 & n872);
  assign n1771 = n1769 & n1770;
  assign n1772 = (n1766 & ~n1768) | (n1766 & n1771) | (~n1768 & n1771);
  assign n1773 = (x132 & x133) | (x132 & ~n1772) | (x133 & ~n1772);
  assign n1774 = n1765 & ~n1773;
  assign n1775 = (x130 & ~x131) | (x130 & n875) | (~x131 & n875);
  assign n1776 = (x130 & x131) | (x130 & ~n877) | (x131 & ~n877);
  assign n1777 = n1775 & n1776;
  assign n1778 = (x130 & x131) | (x130 & n883) | (x131 & n883);
  assign n1779 = (~x130 & x131) | (~x130 & n885) | (x131 & n885);
  assign n1780 = n1778 & n1779;
  assign n1781 = (n1775 & ~n1777) | (n1775 & n1780) | (~n1777 & n1780);
  assign n1782 = (x132 & x133) | (x132 & n1781) | (x133 & n1781);
  assign n1783 = (x130 & ~x131) | (x130 & n888) | (~x131 & n888);
  assign n1784 = (x130 & x131) | (x130 & ~n890) | (x131 & ~n890);
  assign n1785 = n1783 & n1784;
  assign n1786 = (x130 & x131) | (x130 & n895) | (x131 & n895);
  assign n1787 = (~x130 & x131) | (~x130 & n897) | (x131 & n897);
  assign n1788 = n1786 & n1787;
  assign n1789 = (n1783 & ~n1785) | (n1783 & n1788) | (~n1785 & n1788);
  assign n1790 = (~x132 & x133) | (~x132 & n1789) | (x133 & n1789);
  assign n1791 = n1782 & n1790;
  assign n1792 = n1774 | n1791;
  assign n1793 = (x130 & ~x131) | (x130 & n945) | (~x131 & n945);
  assign n1794 = (x130 & x131) | (x130 & ~n947) | (x131 & ~n947);
  assign n1795 = n1793 & n1794;
  assign n1796 = (x130 & x131) | (x130 & n909) | (x131 & n909);
  assign n1797 = (~x130 & x131) | (~x130 & n911) | (x131 & n911);
  assign n1798 = n1796 & n1797;
  assign n1799 = (n1793 & ~n1795) | (n1793 & n1798) | (~n1795 & n1798);
  assign n1800 = (x132 & x133) | (x132 & ~n1799) | (x133 & ~n1799);
  assign n1801 = (x130 & ~x131) | (x130 & n900) | (~x131 & n900);
  assign n1802 = (x130 & x131) | (x130 & ~n902) | (x131 & ~n902);
  assign n1803 = n1801 & n1802;
  assign n1804 = (x130 & x131) | (x130 & n940) | (x131 & n940);
  assign n1805 = (~x130 & x131) | (~x130 & n942) | (x131 & n942);
  assign n1806 = n1804 & n1805;
  assign n1807 = (n1801 & ~n1803) | (n1801 & n1806) | (~n1803 & n1806);
  assign n1808 = (x132 & ~x133) | (x132 & n1807) | (~x133 & n1807);
  assign n1809 = ~n1800 & n1808;
  assign n1810 = (x130 & ~x131) | (x130 & n931) | (~x131 & n931);
  assign n1811 = (x130 & x131) | (x130 & ~n933) | (x131 & ~n933);
  assign n1812 = n1810 & n1811;
  assign n1813 = (x130 & x131) | (x130 & n952) | (x131 & n952);
  assign n1814 = (~x130 & x131) | (~x130 & n954) | (x131 & n954);
  assign n1815 = n1813 & n1814;
  assign n1816 = (n1810 & ~n1812) | (n1810 & n1815) | (~n1812 & n1815);
  assign n1817 = (~x132 & x133) | (~x132 & n1816) | (x133 & n1816);
  assign n1818 = (x130 & ~x131) | (x130 & n917) | (~x131 & n917);
  assign n1819 = (x130 & x131) | (x130 & ~n921) | (x131 & ~n921);
  assign n1820 = n1818 & n1819;
  assign n1821 = (x130 & x131) | (x130 & n926) | (x131 & n926);
  assign n1822 = (~x130 & x131) | (~x130 & n928) | (x131 & n928);
  assign n1823 = n1821 & n1822;
  assign n1824 = (n1818 & ~n1820) | (n1818 & n1823) | (~n1820 & n1823);
  assign n1825 = (x132 & x133) | (x132 & n1824) | (x133 & n1824);
  assign n1826 = n1809 | n1825;
  assign n1827 = (n1809 & n1817) | (n1809 & n1826) | (n1817 & n1826);
  assign n1828 = x134 & ~n1827;
  assign n1829 = x134 & ~n1792;
  assign n1830 = (n1792 & ~n1828) | (n1792 & n1829) | (~n1828 & n1829);
  assign n1831 = (x130 & ~x131) | (x130 & n1218) | (~x131 & n1218);
  assign n1832 = (x130 & x131) | (x130 & ~n1228) | (x131 & ~n1228);
  assign n1833 = n1831 & n1832;
  assign n1834 = (x130 & x131) | (x130 & n1022) | (x131 & n1022);
  assign n1835 = (~x130 & x131) | (~x130 & n1031) | (x131 & n1031);
  assign n1836 = n1834 & n1835;
  assign n1837 = (n1831 & ~n1833) | (n1831 & n1836) | (~n1833 & n1836);
  assign n1838 = (x132 & ~x133) | (x132 & n1837) | (~x133 & n1837);
  assign n1839 = (x130 & ~x131) | (x130 & n1042) | (~x131 & n1042);
  assign n1840 = (x130 & x131) | (x130 & ~n1051) | (x131 & ~n1051);
  assign n1841 = n1839 & n1840;
  assign n1842 = (x130 & x131) | (x130 & n1073) | (x131 & n1073);
  assign n1843 = (~x130 & x131) | (~x130 & n1083) | (x131 & n1083);
  assign n1844 = n1842 & n1843;
  assign n1845 = (n1839 & ~n1841) | (n1839 & n1844) | (~n1841 & n1844);
  assign n1846 = (x132 & x133) | (x132 & ~n1845) | (x133 & ~n1845);
  assign n1847 = n1838 & ~n1846;
  assign n1848 = (x130 & ~x131) | (x130 & n1065) | (~x131 & n1065);
  assign n1849 = (x130 & x131) | (x130 & ~n1094) | (x131 & ~n1094);
  assign n1850 = n1848 & n1849;
  assign n1851 = (x130 & x131) | (x130 & n1117) | (x131 & n1117);
  assign n1852 = (~x130 & x131) | (~x130 & n1127) | (x131 & n1127);
  assign n1853 = n1851 & n1852;
  assign n1854 = (n1848 & ~n1850) | (n1848 & n1853) | (~n1850 & n1853);
  assign n1855 = (x132 & x133) | (x132 & n1854) | (x133 & n1854);
  assign n1856 = (x130 & ~x131) | (x130 & n1107) | (~x131 & n1107);
  assign n1857 = (x130 & x131) | (x130 & ~n1137) | (x131 & ~n1137);
  assign n1858 = n1856 & n1857;
  assign n1859 = (x130 & x131) | (x130 & n978) | (x131 & n978);
  assign n1860 = (~x130 & x131) | (~x130 & n988) | (x131 & n988);
  assign n1861 = n1859 & n1860;
  assign n1862 = (n1856 & ~n1858) | (n1856 & n1861) | (~n1858 & n1861);
  assign n1863 = (~x132 & x133) | (~x132 & n1862) | (x133 & n1862);
  assign n1864 = n1855 & n1863;
  assign n1865 = n1847 | n1864;
  assign n1866 = (x130 & x131) | (x130 & n1305) | (x131 & n1305);
  assign n1867 = (x130 & x131) | (x130 & ~n1242) | (x131 & ~n1242);
  assign n1868 = n1553 & ~n1867;
  assign n1869 = n1565 | n1868;
  assign n1870 = (n1866 & n1868) | (n1866 & n1869) | (n1868 & n1869);
  assign n1871 = (x132 & x133) | (x132 & ~n1870) | (x133 & ~n1870);
  assign n1872 = (x130 & ~x131) | (x130 & n999) | (~x131 & n999);
  assign n1873 = (x130 & x131) | (x130 & ~n1009) | (x131 & ~n1009);
  assign n1874 = n1872 & n1873;
  assign n1875 = (x130 & x131) | (x130 & n1275) | (x131 & n1275);
  assign n1876 = (~x130 & x131) | (~x130 & n1284) | (x131 & n1284);
  assign n1877 = n1875 & n1876;
  assign n1878 = (n1872 & ~n1874) | (n1872 & n1877) | (~n1874 & n1877);
  assign n1879 = (x132 & ~x133) | (x132 & n1878) | (~x133 & n1878);
  assign n1880 = ~n1871 & n1879;
  assign n1881 = (x130 & ~x131) | (x130 & n1174) | (~x131 & n1174);
  assign n1882 = (x130 & x131) | (x130 & ~n1184) | (x131 & ~n1184);
  assign n1883 = n1881 & n1882;
  assign n1884 = (x130 & x131) | (x130 & n1197) | (x131 & n1197);
  assign n1885 = (~x130 & x131) | (~x130 & n1207) | (x131 & n1207);
  assign n1886 = n1884 & n1885;
  assign n1887 = (n1881 & ~n1883) | (n1881 & n1886) | (~n1883 & n1886);
  assign n1888 = (~x132 & x133) | (~x132 & n1887) | (x133 & n1887);
  assign n1889 = (x130 & x131) | (x130 & ~n1262) | (x131 & ~n1262);
  assign n1890 = n1562 & n1889;
  assign n1891 = (x130 & x131) | (x130 & n1153) | (x131 & n1153);
  assign n1892 = (~x130 & x131) | (~x130 & n1163) | (x131 & n1163);
  assign n1893 = n1891 & n1892;
  assign n1894 = (n1562 & ~n1890) | (n1562 & n1893) | (~n1890 & n1893);
  assign n1895 = (x132 & x133) | (x132 & n1894) | (x133 & n1894);
  assign n1896 = n1880 | n1895;
  assign n1897 = (n1880 & n1888) | (n1880 & n1896) | (n1888 & n1896);
  assign n1898 = x134 & ~n1897;
  assign n1899 = x134 & ~n1865;
  assign n1900 = (n1865 & ~n1898) | (n1865 & n1899) | (~n1898 & n1899);
  assign n1901 = (x130 & x131) | (x130 & n219) | (x131 & n219);
  assign n1902 = (~x130 & x131) | (~x130 & n233) | (x131 & n233);
  assign n1903 = n1901 & n1902;
  assign n1904 = x130 & n209;
  assign n1905 = ~x130 & n198;
  assign n1906 = (~x131 & n1904) | (~x131 & n1905) | (n1904 & n1905);
  assign n1907 = n1903 | n1906;
  assign n1908 = (x132 & x133) | (x132 & n1907) | (x133 & n1907);
  assign n1909 = (x130 & x131) | (x130 & n264) | (x131 & n264);
  assign n1910 = (~x130 & x131) | (~x130 & n277) | (x131 & n277);
  assign n1911 = n1909 & n1910;
  assign n1912 = x130 & n254;
  assign n1913 = ~x130 & n243;
  assign n1914 = (~x131 & n1912) | (~x131 & n1913) | (n1912 & n1913);
  assign n1915 = n1911 | n1914;
  assign n1916 = (~x132 & x133) | (~x132 & n1915) | (x133 & n1915);
  assign n1917 = n1908 & n1916;
  assign n1918 = (x130 & x131) | (x130 & n175) | (x131 & n175);
  assign n1919 = (~x130 & x131) | (~x130 & n188) | (x131 & n188);
  assign n1920 = n1918 & n1919;
  assign n1921 = x130 & n165;
  assign n1922 = ~x130 & n154;
  assign n1923 = (~x131 & n1921) | (~x131 & n1922) | (n1921 & n1922);
  assign n1924 = n1920 | n1923;
  assign n1925 = x132 & n1924;
  assign n1926 = (x131 & n1379) | (x131 & n1380) | (n1379 & n1380);
  assign n1927 = (x130 & x131) | (x130 & ~n479) | (x131 & ~n479);
  assign n1928 = (x130 & ~x131) | (x130 & n468) | (~x131 & n468);
  assign n1929 = n1926 | n1928;
  assign n1930 = (n1926 & ~n1927) | (n1926 & n1929) | (~n1927 & n1929);
  assign n1931 = ~x132 & n1930;
  assign n1932 = (~x133 & n1925) | (~x133 & n1931) | (n1925 & n1931);
  assign n1933 = n1917 | n1932;
  assign n1934 = (x131 & n1318) | (x131 & n1319) | (n1318 & n1319);
  assign n1935 = (x130 & x131) | (x130 & ~n390) | (x131 & ~n390);
  assign n1936 = (x130 & ~x131) | (x130 & n379) | (~x131 & n379);
  assign n1937 = n1934 | n1936;
  assign n1938 = (n1934 & ~n1935) | (n1934 & n1937) | (~n1935 & n1937);
  assign n1939 = (x132 & x133) | (x132 & ~n1938) | (x133 & ~n1938);
  assign n1940 = (x130 & x131) | (x130 & n308) | (x131 & n308);
  assign n1941 = (~x130 & x131) | (~x130 & n369) | (x131 & n369);
  assign n1942 = n1940 & n1941;
  assign n1943 = x130 & n298;
  assign n1944 = ~x130 & n287;
  assign n1945 = (~x131 & n1943) | (~x131 & n1944) | (n1943 & n1944);
  assign n1946 = n1942 | n1945;
  assign n1947 = (x132 & ~x133) | (x132 & n1946) | (~x133 & n1946);
  assign n1948 = ~n1939 & n1947;
  assign n1949 = (x130 & x131) | (x130 & n446) | (x131 & n446);
  assign n1950 = (~x130 & x131) | (~x130 & n458) | (x131 & n458);
  assign n1951 = n1949 & ~n1950;
  assign n1952 = x130 & n436;
  assign n1953 = ~x130 & n425;
  assign n1954 = (~x131 & n1952) | (~x131 & n1953) | (n1952 & n1953);
  assign n1955 = (n1949 & ~n1951) | (n1949 & n1954) | (~n1951 & n1954);
  assign n1956 = (~x132 & x133) | (~x132 & n1955) | (x133 & n1955);
  assign n1957 = (x130 & x131) | (x130 & n356) | (x131 & n356);
  assign n1958 = (~x130 & x131) | (~x130 & n415) | (x131 & n415);
  assign n1959 = n1957 & n1958;
  assign n1960 = x130 & n346;
  assign n1961 = ~x130 & n333;
  assign n1962 = (~x131 & n1960) | (~x131 & n1961) | (n1960 & n1961);
  assign n1963 = n1959 | n1962;
  assign n1964 = (x132 & x133) | (x132 & n1963) | (x133 & n1963);
  assign n1965 = n1948 | n1964;
  assign n1966 = (n1948 & n1956) | (n1948 & n1965) | (n1956 & n1965);
  assign n1967 = x134 & ~n1966;
  assign n1968 = x134 & ~n1933;
  assign n1969 = (n1933 & ~n1967) | (n1933 & n1968) | (~n1967 & n1968);
  assign n1970 = (x130 & x131) | (x130 & n582) | (x131 & n582);
  assign n1971 = (~x130 & x131) | (~x130 & n596) | (x131 & n596);
  assign n1972 = n1970 & n1971;
  assign n1973 = x130 & n572;
  assign n1974 = ~x130 & n561;
  assign n1975 = (~x131 & n1973) | (~x131 & n1974) | (n1973 & n1974);
  assign n1976 = n1972 | n1975;
  assign n1977 = (x132 & x133) | (x132 & n1976) | (x133 & n1976);
  assign n1978 = (x130 & x131) | (x130 & n627) | (x131 & n627);
  assign n1979 = (~x130 & x131) | (~x130 & n640) | (x131 & n640);
  assign n1980 = n1978 & n1979;
  assign n1981 = x130 & n617;
  assign n1982 = ~x130 & n606;
  assign n1983 = (~x131 & n1981) | (~x131 & n1982) | (n1981 & n1982);
  assign n1984 = n1980 | n1983;
  assign n1985 = (~x132 & x133) | (~x132 & n1984) | (x133 & n1984);
  assign n1986 = n1977 & n1985;
  assign n1987 = (x130 & x131) | (x130 & n538) | (x131 & n538);
  assign n1988 = (~x130 & x131) | (~x130 & n551) | (x131 & n551);
  assign n1989 = n1987 & n1988;
  assign n1990 = x130 & n528;
  assign n1991 = ~x130 & n517;
  assign n1992 = (~x131 & n1990) | (~x131 & n1991) | (n1990 & n1991);
  assign n1993 = n1989 | n1992;
  assign n1994 = x132 & n1993;
  assign n1995 = (x131 & n1452) | (x131 & n1453) | (n1452 & n1453);
  assign n1996 = (x130 & x131) | (x130 & ~n837) | (x131 & ~n837);
  assign n1997 = (x130 & ~x131) | (x130 & n826) | (~x131 & n826);
  assign n1998 = n1995 | n1997;
  assign n1999 = (n1995 & ~n1996) | (n1995 & n1998) | (~n1996 & n1998);
  assign n2000 = ~x132 & n1999;
  assign n2001 = (~x133 & n1994) | (~x133 & n2000) | (n1994 & n2000);
  assign n2002 = n1986 | n2001;
  assign n2003 = (x131 & n1391) | (x131 & n1392) | (n1391 & n1392);
  assign n2004 = (x130 & x131) | (x130 & ~n793) | (x131 & ~n793);
  assign n2005 = (x130 & ~x131) | (x130 & n782) | (~x131 & n782);
  assign n2006 = n2003 | n2005;
  assign n2007 = (n2003 & ~n2004) | (n2003 & n2006) | (~n2004 & n2006);
  assign n2008 = (x132 & x133) | (x132 & ~n2007) | (x133 & ~n2007);
  assign n2009 = (x130 & x131) | (x130 & n671) | (x131 & n671);
  assign n2010 = (~x130 & x131) | (~x130 & n772) | (x131 & n772);
  assign n2011 = n2009 & n2010;
  assign n2012 = x130 & n661;
  assign n2013 = ~x130 & n650;
  assign n2014 = (~x131 & n2012) | (~x131 & n2013) | (n2012 & n2013);
  assign n2015 = n2011 | n2014;
  assign n2016 = (x132 & ~x133) | (x132 & n2015) | (~x133 & n2015);
  assign n2017 = ~n2008 & n2016;
  assign n2018 = (x130 & x131) | (x130 & n756) | (x131 & n756);
  assign n2019 = (~x130 & x131) | (~x130 & n816) | (x131 & n816);
  assign n2020 = n2018 & ~n2019;
  assign n2021 = x130 & n746;
  assign n2022 = ~x130 & n735;
  assign n2023 = (~x131 & n2021) | (~x131 & n2022) | (n2021 & n2022);
  assign n2024 = (n2018 & ~n2020) | (n2018 & n2023) | (~n2020 & n2023);
  assign n2025 = (~x132 & x133) | (~x132 & n2024) | (x133 & n2024);
  assign n2026 = (x130 & x131) | (x130 & n712) | (x131 & n712);
  assign n2027 = (~x130 & x131) | (~x130 & n725) | (x131 & n725);
  assign n2028 = n2026 & n2027;
  assign n2029 = (x130 & x131) | (x130 & ~n702) | (x131 & ~n702);
  assign n2030 = (x130 & ~x131) | (x130 & n693) | (~x131 & n693);
  assign n2031 = n2029 | n2030;
  assign n2032 = (n2028 & ~n2029) | (n2028 & n2031) | (~n2029 & n2031);
  assign n2033 = (x132 & x133) | (x132 & n2032) | (x133 & n2032);
  assign n2034 = n2017 | n2033;
  assign n2035 = (n2017 & n2025) | (n2017 & n2034) | (n2025 & n2034);
  assign n2036 = x134 & ~n2035;
  assign n2037 = x134 & ~n2002;
  assign n2038 = (n2002 & ~n2036) | (n2002 & n2037) | (~n2036 & n2037);
  assign n2039 = (x130 & x131) | (x130 & n877) | (x131 & n877);
  assign n2040 = (~x130 & x131) | (~x130 & n883) | (x131 & n883);
  assign n2041 = n2039 & n2040;
  assign n2042 = x130 & n875;
  assign n2043 = ~x130 & n872;
  assign n2044 = (~x131 & n2042) | (~x131 & n2043) | (n2042 & n2043);
  assign n2045 = n2041 | n2044;
  assign n2046 = (x132 & x133) | (x132 & n2045) | (x133 & n2045);
  assign n2047 = (x130 & x131) | (x130 & n890) | (x131 & n890);
  assign n2048 = (~x130 & x131) | (~x130 & n895) | (x131 & n895);
  assign n2049 = n2047 & n2048;
  assign n2050 = x130 & n888;
  assign n2051 = ~x130 & n885;
  assign n2052 = (~x131 & n2050) | (~x131 & n2051) | (n2050 & n2051);
  assign n2053 = n2049 | n2052;
  assign n2054 = (~x132 & x133) | (~x132 & n2053) | (x133 & n2053);
  assign n2055 = n2046 & n2054;
  assign n2056 = (x130 & x131) | (x130 & n865) | (x131 & n865);
  assign n2057 = (~x130 & x131) | (~x130 & n870) | (x131 & n870);
  assign n2058 = n2056 & n2057;
  assign n2059 = x130 & n863;
  assign n2060 = ~x130 & n860;
  assign n2061 = (~x131 & n2059) | (~x131 & n2060) | (n2059 & n2060);
  assign n2062 = n2058 | n2061;
  assign n2063 = x132 & n2062;
  assign n2064 = (x131 & n1525) | (x131 & n1526) | (n1525 & n1526);
  assign n2065 = (x130 & x131) | (x130 & ~n957) | (x131 & ~n957);
  assign n2066 = (x130 & ~x131) | (x130 & n954) | (~x131 & n954);
  assign n2067 = n2064 | n2066;
  assign n2068 = (n2064 & ~n2065) | (n2064 & n2067) | (~n2065 & n2067);
  assign n2069 = ~x132 & n2068;
  assign n2070 = (~x133 & n2063) | (~x133 & n2069) | (n2063 & n2069);
  assign n2071 = n2055 | n2070;
  assign n2072 = (x131 & n1464) | (x131 & n1465) | (n1464 & n1465);
  assign n2073 = (x130 & x131) | (x130 & ~n945) | (x131 & ~n945);
  assign n2074 = (x130 & ~x131) | (x130 & n942) | (~x131 & n942);
  assign n2075 = n2072 | n2074;
  assign n2076 = (n2072 & ~n2073) | (n2072 & n2075) | (~n2073 & n2075);
  assign n2077 = (x132 & x133) | (x132 & ~n2076) | (x133 & ~n2076);
  assign n2078 = (x130 & x131) | (x130 & n902) | (x131 & n902);
  assign n2079 = (~x130 & x131) | (~x130 & n940) | (x131 & n940);
  assign n2080 = n2078 & n2079;
  assign n2081 = x130 & n900;
  assign n2082 = ~x130 & n897;
  assign n2083 = (~x131 & n2081) | (~x131 & n2082) | (n2081 & n2082);
  assign n2084 = n2080 | n2083;
  assign n2085 = (x132 & ~x133) | (x132 & n2084) | (~x133 & n2084);
  assign n2086 = ~n2077 & n2085;
  assign n2087 = (x130 & x131) | (x130 & n933) | (x131 & n933);
  assign n2088 = (~x130 & x131) | (~x130 & n952) | (x131 & n952);
  assign n2089 = n2087 & ~n2088;
  assign n2090 = x130 & n931;
  assign n2091 = ~x130 & n928;
  assign n2092 = (~x131 & n2090) | (~x131 & n2091) | (n2090 & n2091);
  assign n2093 = (n2087 & ~n2089) | (n2087 & n2092) | (~n2089 & n2092);
  assign n2094 = (~x132 & x133) | (~x132 & n2093) | (x133 & n2093);
  assign n2095 = (x130 & x131) | (x130 & n921) | (x131 & n921);
  assign n2096 = (~x130 & x131) | (~x130 & n926) | (x131 & n926);
  assign n2097 = n2095 & n2096;
  assign n2098 = x130 & n917;
  assign n2099 = ~x130 & n911;
  assign n2100 = (~x131 & n2098) | (~x131 & n2099) | (n2098 & n2099);
  assign n2101 = n2097 | n2100;
  assign n2102 = (x132 & x133) | (x132 & n2101) | (x133 & n2101);
  assign n2103 = n2086 | n2102;
  assign n2104 = (n2086 & n2094) | (n2086 & n2103) | (n2094 & n2103);
  assign n2105 = x134 & ~n2104;
  assign n2106 = x134 & ~n2071;
  assign n2107 = (n2071 & ~n2105) | (n2071 & n2106) | (~n2105 & n2106);
  assign n2108 = (x130 & x131) | (x130 & n1094) | (x131 & n1094);
  assign n2109 = (~x130 & x131) | (~x130 & n1117) | (x131 & n1117);
  assign n2110 = n2108 & n2109;
  assign n2111 = x130 & n1065;
  assign n2112 = ~x130 & n1083;
  assign n2113 = (~x131 & n2111) | (~x131 & n2112) | (n2111 & n2112);
  assign n2114 = n2110 | n2113;
  assign n2115 = (x132 & x133) | (x132 & n2114) | (x133 & n2114);
  assign n2116 = (x131 & n1593) | (x131 & n1594) | (n1593 & n1594);
  assign n2117 = (x130 & x131) | (x130 & ~n1107) | (x131 & ~n1107);
  assign n2118 = (x130 & ~x131) | (x130 & n1127) | (~x131 & n1127);
  assign n2119 = n2116 | n2118;
  assign n2120 = (n2116 & ~n2117) | (n2116 & n2119) | (~n2117 & n2119);
  assign n2121 = (~x132 & x133) | (~x132 & n2120) | (x133 & n2120);
  assign n2122 = n2115 & n2121;
  assign n2123 = (x130 & x131) | (x130 & n1051) | (x131 & n1051);
  assign n2124 = (~x130 & x131) | (~x130 & n1073) | (x131 & n1073);
  assign n2125 = n2123 & n2124;
  assign n2126 = x130 & n1042;
  assign n2127 = ~x130 & n1031;
  assign n2128 = (~x131 & n2126) | (~x131 & n2127) | (n2126 & n2127);
  assign n2129 = n2125 | n2128;
  assign n2130 = x132 & n2129;
  assign n2131 = (x131 & n1584) | (x131 & n1585) | (n1584 & n1585);
  assign n2132 = (x130 & x131) | (x130 & ~n1218) | (x131 & ~n1218);
  assign n2133 = (x130 & ~x131) | (x130 & n1207) | (~x131 & n1207);
  assign n2134 = n2131 | n2133;
  assign n2135 = (n2131 & ~n2132) | (n2131 & n2134) | (~n2132 & n2134);
  assign n2136 = ~x132 & n2135;
  assign n2137 = (~x133 & n2130) | (~x133 & n2136) | (n2130 & n2136);
  assign n2138 = n2122 | n2137;
  assign n2139 = x130 & n1242;
  assign n2140 = (x131 & n1560) | (x131 & n2139) | (n1560 & n2139);
  assign n2141 = x131 & ~n2140;
  assign n2142 = (~x130 & n1284) | (~x130 & n1296) | (n1284 & n1296);
  assign n2143 = (~x131 & n1296) | (~x131 & n2142) | (n1296 & n2142);
  assign n2144 = (n2140 & ~n2141) | (n2140 & n2143) | (~n2141 & n2143);
  assign n2145 = (x132 & x133) | (x132 & ~n2144) | (x133 & ~n2144);
  assign n2146 = (x130 & x131) | (x130 & n1009) | (x131 & n1009);
  assign n2147 = (~x130 & x131) | (~x130 & n1275) | (x131 & n1275);
  assign n2148 = n2146 & n2147;
  assign n2149 = x130 & n999;
  assign n2150 = ~x130 & n988;
  assign n2151 = (~x131 & n2149) | (~x131 & n2150) | (n2149 & n2150);
  assign n2152 = n2148 | n2151;
  assign n2153 = (x132 & ~x133) | (x132 & n2152) | (~x133 & n2152);
  assign n2154 = ~n2145 & n2153;
  assign n2155 = (x130 & x131) | (x130 & n1184) | (x131 & n1184);
  assign n2156 = (~x130 & x131) | (~x130 & n1197) | (x131 & n1197);
  assign n2157 = n2155 & ~n2156;
  assign n2158 = x130 & n1174;
  assign n2159 = ~x130 & n1163;
  assign n2160 = (~x131 & n2158) | (~x131 & n2159) | (n2158 & n2159);
  assign n2161 = (n2155 & ~n2157) | (n2155 & n2160) | (~n2157 & n2160);
  assign n2162 = (~x132 & x133) | (~x132 & n2161) | (x133 & n2161);
  assign n2163 = (x131 & n1537) | (x131 & n1538) | (n1537 & n1538);
  assign n2164 = (x130 & x131) | (x130 & ~n1253) | (x131 & ~n1253);
  assign n2165 = n1565 | n2163;
  assign n2166 = (n2163 & ~n2164) | (n2163 & n2165) | (~n2164 & n2165);
  assign n2167 = (x132 & x133) | (x132 & n2166) | (x133 & n2166);
  assign n2168 = n2154 | n2167;
  assign n2169 = (n2154 & n2162) | (n2154 & n2168) | (n2162 & n2168);
  assign n2170 = x134 & ~n2169;
  assign n2171 = x134 & ~n2138;
  assign n2172 = (n2138 & ~n2170) | (n2138 & n2171) | (~n2170 & n2171);
  assign n2173 = x133 | n403;
  assign n2174 = (x132 & ~x133) | (x132 & n359) | (~x133 & n359);
  assign n2175 = n359 & ~n2174;
  assign n2176 = (n678 & n2173) | (n678 & n2175) | (n2173 & n2175);
  assign n2177 = x133 | n311;
  assign n2178 = (x132 & x133) | (x132 & ~n449) | (x133 & ~n449);
  assign n2179 = n449 & n2178;
  assign n2180 = (~n763 & n2177) | (~n763 & n2179) | (n2177 & n2179);
  assign n2181 = n2176 | n2180;
  assign n2182 = x134 & ~n2181;
  assign n2183 = (x132 & x133) | (x132 & ~n178) | (x133 & ~n178);
  assign n2184 = n493 & ~n2183;
  assign n2185 = x133 | n2184;
  assign n2186 = (x132 & ~x133) | (x132 & n267) | (~x133 & n267);
  assign n2187 = (~x132 & n222) | (~x132 & n2186) | (n222 & n2186);
  assign n2188 = (n2184 & n2185) | (n2184 & n2186) | (n2185 & n2186);
  assign n2189 = (n2185 & n2187) | (n2185 & n2188) | (n2187 & n2188);
  assign n2190 = x134 & ~n2189;
  assign n2191 = (~n2182 & n2189) | (~n2182 & n2190) | (n2189 & n2190);
  assign n2192 = (x132 & x133) | (x132 & ~n806) | (x133 & ~n806);
  assign n2193 = (x132 & ~x133) | (x132 & n674) | (~x133 & n674);
  assign n2194 = ~n2192 & n2193;
  assign n2195 = (~x132 & x133) | (~x132 & n759) | (x133 & n759);
  assign n2196 = (x132 & x133) | (x132 & n715) | (x133 & n715);
  assign n2197 = n2194 | n2196;
  assign n2198 = (n2194 & n2195) | (n2194 & n2197) | (n2195 & n2197);
  assign n2199 = x134 & ~n2198;
  assign n2200 = (~x132 & x133) | (~x132 & n630) | (x133 & n630);
  assign n2201 = x132 & n541;
  assign n2202 = ~x132 & n850;
  assign n2203 = (~x133 & n2201) | (~x133 & n2202) | (n2201 & n2202);
  assign n2204 = (x132 & x133) | (x132 & n585) | (x133 & n585);
  assign n2205 = n2203 | n2204;
  assign n2206 = (n2200 & n2203) | (n2200 & n2205) | (n2203 & n2205);
  assign n2207 = x134 & ~n2206;
  assign n2208 = (~n2199 & n2206) | (~n2199 & n2207) | (n2206 & n2207);
  assign n2209 = (x132 & x133) | (x132 & ~n950) | (x133 & ~n950);
  assign n2210 = (x132 & ~x133) | (x132 & n905) | (~x133 & n905);
  assign n2211 = ~n2209 & n2210;
  assign n2212 = (~x132 & x133) | (~x132 & n936) | (x133 & n936);
  assign n2213 = (x132 & x133) | (x132 & n924) | (x133 & n924);
  assign n2214 = n2211 | n2213;
  assign n2215 = (n2211 & n2212) | (n2211 & n2214) | (n2212 & n2214);
  assign n2216 = x134 & ~n2215;
  assign n2217 = (~x132 & x133) | (~x132 & n893) | (x133 & n893);
  assign n2218 = x132 & n868;
  assign n2219 = ~x132 & n962;
  assign n2220 = (~x133 & n2218) | (~x133 & n2219) | (n2218 & n2219);
  assign n2221 = (x132 & x133) | (x132 & n880) | (x133 & n880);
  assign n2222 = n2220 | n2221;
  assign n2223 = (n2217 & n2220) | (n2217 & n2222) | (n2220 & n2222);
  assign n2224 = x134 & ~n2223;
  assign n2225 = (~n2216 & n2223) | (~n2216 & n2224) | (n2223 & n2224);
  assign n2226 = (x132 & x133) | (x132 & ~n1310) | (x133 & ~n1310);
  assign n2227 = n1013 & ~n2226;
  assign n2228 = (~x132 & x133) | (~x132 & n1187) | (x133 & n1187);
  assign n2229 = (x132 & x133) | (x132 & n1265) | (x133 & n1265);
  assign n2230 = n2227 | n2229;
  assign n2231 = (n2227 & n2228) | (n2227 & n2230) | (n2228 & n2230);
  assign n2232 = x134 & ~n2231;
  assign n2233 = (x132 & x133) | (x132 & n1097) | (x133 & n1097);
  assign n2234 = (~x132 & x133) | (~x132 & n1140) | (x133 & n1140);
  assign n2235 = n2233 & n2234;
  assign n2236 = (x132 & ~x133) | (x132 & n1231) | (~x133 & n1231);
  assign n2237 = (x132 & x133) | (x132 & ~n1054) | (x133 & ~n1054);
  assign n2238 = ~n2235 & n2237;
  assign n2239 = (n2235 & n2236) | (n2235 & ~n2238) | (n2236 & ~n2238);
  assign n2240 = x134 & ~n2239;
  assign n2241 = (~n2232 & n2239) | (~n2232 & n2240) | (n2239 & n2240);
  assign n2242 = (x132 & ~x133) | (x132 & n1340) | (~x133 & n1340);
  assign n2243 = (x132 & x133) | (x132 & ~n1384) | (x133 & ~n1384);
  assign n2244 = n2242 & ~n2243;
  assign n2245 = (x132 & x133) | (x132 & n1376) | (x133 & n1376);
  assign n2246 = (~x132 & x133) | (~x132 & n1359) | (x133 & n1359);
  assign n2247 = n2245 & n2246;
  assign n2248 = n2244 | n2247;
  assign n2249 = ~n1324 & n1368;
  assign n2250 = (x132 & ~x133) | (x132 & n1348) | (~x133 & n1348);
  assign n2251 = (x132 & x133) | (x132 & n1331) | (x133 & n1331);
  assign n2252 = (n2249 & n2250) | (n2249 & n2251) | (n2250 & n2251);
  assign n2253 = n2249 | n2252;
  assign n2254 = x134 & ~n2253;
  assign n2255 = x134 & ~n2248;
  assign n2256 = (n2248 & ~n2254) | (n2248 & n2255) | (~n2254 & n2255);
  assign n2257 = (x132 & ~x133) | (x132 & n1413) | (~x133 & n1413);
  assign n2258 = (x132 & x133) | (x132 & ~n1457) | (x133 & ~n1457);
  assign n2259 = n2257 & ~n2258;
  assign n2260 = (x132 & x133) | (x132 & n1449) | (x133 & n1449);
  assign n2261 = (~x132 & x133) | (~x132 & n1432) | (x133 & n1432);
  assign n2262 = n2260 & n2261;
  assign n2263 = n2259 | n2262;
  assign n2264 = ~n1397 & n1441;
  assign n2265 = (x132 & ~x133) | (x132 & n1421) | (~x133 & n1421);
  assign n2266 = (x132 & x133) | (x132 & n1404) | (x133 & n1404);
  assign n2267 = (n2264 & n2265) | (n2264 & n2266) | (n2265 & n2266);
  assign n2268 = n2264 | n2267;
  assign n2269 = x134 & ~n2268;
  assign n2270 = x134 & ~n2263;
  assign n2271 = (n2263 & ~n2269) | (n2263 & n2270) | (~n2269 & n2270);
  assign n2272 = (x132 & ~x133) | (x132 & n1486) | (~x133 & n1486);
  assign n2273 = (x132 & x133) | (x132 & ~n1530) | (x133 & ~n1530);
  assign n2274 = n2272 & ~n2273;
  assign n2275 = (x132 & x133) | (x132 & n1522) | (x133 & n1522);
  assign n2276 = (~x132 & x133) | (~x132 & n1505) | (x133 & n1505);
  assign n2277 = n2275 & n2276;
  assign n2278 = n2274 | n2277;
  assign n2279 = ~n1470 & n1514;
  assign n2280 = (x132 & ~x133) | (x132 & n1494) | (~x133 & n1494);
  assign n2281 = (x132 & x133) | (x132 & n1477) | (x133 & n1477);
  assign n2282 = (n2279 & n2280) | (n2279 & n2281) | (n2280 & n2281);
  assign n2283 = n2279 | n2282;
  assign n2284 = x134 & ~n2283;
  assign n2285 = x134 & ~n2278;
  assign n2286 = (n2278 & ~n2284) | (n2278 & n2285) | (~n2284 & n2285);
  assign n2287 = x133 | n1589;
  assign n2288 = (x132 & ~x133) | (x132 & n1581) | (~x133 & n1581);
  assign n2289 = n1581 & ~n2288;
  assign n2290 = (n678 & n2287) | (n678 & n2289) | (n2287 & n2289);
  assign n2291 = x133 | n1550;
  assign n2292 = (x132 & x133) | (x132 & ~n1606) | (x133 & ~n1606);
  assign n2293 = n1606 & n2292;
  assign n2294 = (~n763 & n2291) | (~n763 & n2293) | (n2291 & n2293);
  assign n2295 = n2290 | n2294;
  assign n2296 = (x132 & ~x133) | (x132 & n1542) | (~x133 & n1542);
  assign n2297 = x133 & n2296;
  assign n2298 = x133 | n1598;
  assign n2299 = (~n763 & n2297) | (~n763 & n2298) | (n2297 & n2298);
  assign n2300 = x133 | n1558;
  assign n2301 = x133 & ~n1571;
  assign n2302 = (n678 & n2300) | (n678 & n2301) | (n2300 & n2301);
  assign n2303 = n2299 | n2302;
  assign n2304 = x134 & ~n2303;
  assign n2305 = x134 & ~n2295;
  assign n2306 = (n2295 & ~n2304) | (n2295 & n2305) | (~n2304 & n2305);
  assign n2307 = x133 | n1662;
  assign n2308 = (x132 & ~x133) | (x132 & n1654) | (~x133 & n1654);
  assign n2309 = n1654 & ~n2308;
  assign n2310 = (n678 & n2307) | (n678 & n2309) | (n2307 & n2309);
  assign n2311 = x133 | n1626;
  assign n2312 = (x132 & x133) | (x132 & ~n1679) | (x133 & ~n1679);
  assign n2313 = n1679 & n2312;
  assign n2314 = (~n763 & n2311) | (~n763 & n2313) | (n2311 & n2313);
  assign n2315 = n2310 | n2314;
  assign n2316 = x133 | n1671;
  assign n2317 = (x132 & ~x133) | (x132 & n1618) | (~x133 & n1618);
  assign n2318 = x133 & n2317;
  assign n2319 = (~n763 & n2316) | (~n763 & n2318) | (n2316 & n2318);
  assign n2320 = x133 | n1635;
  assign n2321 = x133 & ~n1644;
  assign n2322 = (n678 & n2320) | (n678 & n2321) | (n2320 & n2321);
  assign n2323 = n2319 | n2322;
  assign n2324 = x134 & ~n2323;
  assign n2325 = x134 & ~n2315;
  assign n2326 = (n2315 & ~n2324) | (n2315 & n2325) | (~n2324 & n2325);
  assign n2327 = x133 | n1735;
  assign n2328 = (x132 & ~x133) | (x132 & n1727) | (~x133 & n1727);
  assign n2329 = n1727 & ~n2328;
  assign n2330 = (n678 & n2327) | (n678 & n2329) | (n2327 & n2329);
  assign n2331 = x133 | n1699;
  assign n2332 = (x132 & x133) | (x132 & ~n1752) | (x133 & ~n1752);
  assign n2333 = n1752 & n2332;
  assign n2334 = (~n763 & n2331) | (~n763 & n2333) | (n2331 & n2333);
  assign n2335 = n2330 | n2334;
  assign n2336 = x133 | n1744;
  assign n2337 = (x132 & ~x133) | (x132 & n1691) | (~x133 & n1691);
  assign n2338 = x133 & n2337;
  assign n2339 = (~n763 & n2336) | (~n763 & n2338) | (n2336 & n2338);
  assign n2340 = x133 | n1708;
  assign n2341 = x133 & ~n1717;
  assign n2342 = (n678 & n2340) | (n678 & n2341) | (n2340 & n2341);
  assign n2343 = n2339 | n2342;
  assign n2344 = x134 & ~n2343;
  assign n2345 = x134 & ~n2335;
  assign n2346 = (n2335 & ~n2344) | (n2335 & n2345) | (~n2344 & n2345);
  assign n2347 = (x132 & x133) | (x132 & n1772) | (x133 & n1772);
  assign n2348 = (~x132 & x133) | (~x132 & n1781) | (x133 & n1781);
  assign n2349 = n2347 & n2348;
  assign n2350 = x132 & n1764;
  assign n2351 = ~x132 & n1816;
  assign n2352 = (~x133 & n2350) | (~x133 & n2351) | (n2350 & n2351);
  assign n2353 = n2349 | n2352;
  assign n2354 = x133 | n1789;
  assign n2355 = (x132 & ~x133) | (x132 & n1824) | (~x133 & n1824);
  assign n2356 = x133 & n2355;
  assign n2357 = (~n763 & n2354) | (~n763 & n2356) | (n2354 & n2356);
  assign n2358 = x133 | n1807;
  assign n2359 = x133 & ~n1800;
  assign n2360 = (n678 & n2358) | (n678 & n2359) | (n2358 & n2359);
  assign n2361 = n2357 | n2360;
  assign n2362 = x134 & ~n2361;
  assign n2363 = x134 & ~n2353;
  assign n2364 = (n2353 & ~n2362) | (n2353 & n2363) | (~n2362 & n2363);
  assign n2365 = (x132 & x133) | (x132 & n1845) | (x133 & n1845);
  assign n2366 = (~x132 & x133) | (~x132 & n1854) | (x133 & n1854);
  assign n2367 = n2365 & n2366;
  assign n2368 = x132 & n1837;
  assign n2369 = ~x132 & n1887;
  assign n2370 = (~x133 & n2368) | (~x133 & n2369) | (n2368 & n2369);
  assign n2371 = n2367 | n2370;
  assign n2372 = x133 | n1862;
  assign n2373 = (x132 & ~x133) | (x132 & n1894) | (~x133 & n1894);
  assign n2374 = x133 & n2373;
  assign n2375 = (~n763 & n2372) | (~n763 & n2374) | (n2372 & n2374);
  assign n2376 = x133 | n1878;
  assign n2377 = x133 & ~n1871;
  assign n2378 = (n678 & n2376) | (n678 & n2377) | (n2376 & n2377);
  assign n2379 = n2375 | n2378;
  assign n2380 = x134 & ~n2379;
  assign n2381 = x134 & ~n2371;
  assign n2382 = (n2371 & ~n2380) | (n2371 & n2381) | (~n2380 & n2381);
  assign n2383 = (x132 & ~x133) | (x132 & n1955) | (~x133 & n1955);
  assign n2384 = (x132 & x133) | (x132 & ~n1930) | (x133 & ~n1930);
  assign n2385 = n2383 & ~n2384;
  assign n2386 = (x132 & x133) | (x132 & n1924) | (x133 & n1924);
  assign n2387 = (~x132 & x133) | (~x132 & n1907) | (x133 & n1907);
  assign n2388 = n2386 & n2387;
  assign n2389 = n2385 | n2388;
  assign n2390 = x133 | n1915;
  assign n2391 = (x132 & ~x133) | (x132 & n1963) | (~x133 & n1963);
  assign n2392 = x133 & n2391;
  assign n2393 = (~n763 & n2390) | (~n763 & n2392) | (n2390 & n2392);
  assign n2394 = x133 | n1946;
  assign n2395 = x133 & ~n1939;
  assign n2396 = (n678 & n2394) | (n678 & n2395) | (n2394 & n2395);
  assign n2397 = n2393 | n2396;
  assign n2398 = x134 & ~n2397;
  assign n2399 = x134 & ~n2389;
  assign n2400 = (n2389 & ~n2398) | (n2389 & n2399) | (~n2398 & n2399);
  assign n2401 = (x132 & ~x133) | (x132 & n2024) | (~x133 & n2024);
  assign n2402 = (x132 & x133) | (x132 & ~n1999) | (x133 & ~n1999);
  assign n2403 = n2401 & ~n2402;
  assign n2404 = (x132 & x133) | (x132 & n1993) | (x133 & n1993);
  assign n2405 = (~x132 & x133) | (~x132 & n1976) | (x133 & n1976);
  assign n2406 = n2404 & n2405;
  assign n2407 = n2403 | n2406;
  assign n2408 = x133 | n1984;
  assign n2409 = (x132 & ~x133) | (x132 & n2032) | (~x133 & n2032);
  assign n2410 = x133 & n2409;
  assign n2411 = (~n763 & n2408) | (~n763 & n2410) | (n2408 & n2410);
  assign n2412 = x133 | n2015;
  assign n2413 = x133 & ~n2008;
  assign n2414 = (n678 & n2412) | (n678 & n2413) | (n2412 & n2413);
  assign n2415 = n2411 | n2414;
  assign n2416 = x134 & ~n2415;
  assign n2417 = x134 & ~n2407;
  assign n2418 = (n2407 & ~n2416) | (n2407 & n2417) | (~n2416 & n2417);
  assign n2419 = (x132 & ~x133) | (x132 & n2093) | (~x133 & n2093);
  assign n2420 = (x132 & x133) | (x132 & ~n2068) | (x133 & ~n2068);
  assign n2421 = n2419 & ~n2420;
  assign n2422 = (x132 & x133) | (x132 & n2062) | (x133 & n2062);
  assign n2423 = (~x132 & x133) | (~x132 & n2045) | (x133 & n2045);
  assign n2424 = n2422 & n2423;
  assign n2425 = n2421 | n2424;
  assign n2426 = x133 | n2053;
  assign n2427 = (x132 & ~x133) | (x132 & n2101) | (~x133 & n2101);
  assign n2428 = x133 & n2427;
  assign n2429 = (~n763 & n2426) | (~n763 & n2428) | (n2426 & n2428);
  assign n2430 = x133 | n2084;
  assign n2431 = x133 & ~n2077;
  assign n2432 = (n678 & n2430) | (n678 & n2431) | (n2430 & n2431);
  assign n2433 = n2429 | n2432;
  assign n2434 = x134 & ~n2433;
  assign n2435 = x134 & ~n2425;
  assign n2436 = (n2425 & ~n2434) | (n2425 & n2435) | (~n2434 & n2435);
  assign n2437 = (x132 & ~x133) | (x132 & n2161) | (~x133 & n2161);
  assign n2438 = (x132 & x133) | (x132 & ~n2135) | (x133 & ~n2135);
  assign n2439 = n2437 & ~n2438;
  assign n2440 = (x132 & x133) | (x132 & n2129) | (x133 & n2129);
  assign n2441 = (~x132 & x133) | (~x132 & n2114) | (x133 & n2114);
  assign n2442 = n2440 & n2441;
  assign n2443 = n2439 | n2442;
  assign n2444 = (x132 & ~x133) | (x132 & n2166) | (~x133 & n2166);
  assign n2445 = x133 & n2444;
  assign n2446 = x133 | n2120;
  assign n2447 = (~n763 & n2445) | (~n763 & n2446) | (n2445 & n2446);
  assign n2448 = x133 | n2152;
  assign n2449 = x133 & ~n2145;
  assign n2450 = (n678 & n2448) | (n678 & n2449) | (n2448 & n2449);
  assign n2451 = n2447 | n2450;
  assign n2452 = x134 & ~n2451;
  assign n2453 = x134 & ~n2443;
  assign n2454 = (n2443 & ~n2452) | (n2443 & n2453) | (~n2452 & n2453);
  assign n2455 = (x132 & x133) | (x132 & ~n311) | (x133 & ~n311);
  assign n2456 = n2186 & ~n2455;
  assign n2457 = (~x132 & x133) | (~x132 & n359) | (x133 & n359);
  assign n2458 = (x132 & x133) | (x132 & n403) | (x133 & n403);
  assign n2459 = n2456 | n2458;
  assign n2460 = (n2456 & n2457) | (n2456 & n2459) | (n2457 & n2459);
  assign n2461 = x134 & ~n2460;
  assign n2462 = (x132 & x133) | (x132 & ~n492) | (x133 & ~n492);
  assign n2463 = (x132 & ~x133) | (x132 & n449) | (~x133 & n449);
  assign n2464 = n2462 | n2463;
  assign n2465 = (x132 & x133) | (x132 & n178) | (x133 & n178);
  assign n2466 = (~x132 & x133) | (~x132 & n222) | (x133 & n222);
  assign n2467 = n2465 & n2466;
  assign n2468 = (~n2462 & n2464) | (~n2462 & n2467) | (n2464 & n2467);
  assign n2469 = x134 & ~n2468;
  assign n2470 = (~n2461 & n2468) | (~n2461 & n2469) | (n2468 & n2469);
  assign n2471 = x133 | n630;
  assign n2472 = (x132 & ~x133) | (x132 & n715) | (~x133 & n715);
  assign n2473 = x133 & n2472;
  assign n2474 = (~n763 & n2471) | (~n763 & n2473) | (n2471 & n2473);
  assign n2475 = x133 | n674;
  assign n2476 = x133 & ~n2192;
  assign n2477 = (n678 & n2475) | (n678 & n2476) | (n2475 & n2476);
  assign n2478 = n2474 | n2477;
  assign n2479 = x134 & ~n2478;
  assign n2480 = n760 & ~n851;
  assign n2481 = (~x132 & x133) | (~x132 & n585) | (x133 & n585);
  assign n2482 = (x132 & x133) | (x132 & n541) | (x133 & n541);
  assign n2483 = n2480 | n2482;
  assign n2484 = (n2480 & n2481) | (n2480 & n2483) | (n2481 & n2483);
  assign n2485 = x134 & ~n2484;
  assign n2486 = (~n2479 & n2484) | (~n2479 & n2485) | (n2484 & n2485);
  assign n2487 = x133 | n893;
  assign n2488 = (x132 & ~x133) | (x132 & n924) | (~x133 & n924);
  assign n2489 = x133 & n2488;
  assign n2490 = (~n763 & n2487) | (~n763 & n2489) | (n2487 & n2489);
  assign n2491 = x133 | n905;
  assign n2492 = x133 & ~n2209;
  assign n2493 = (n678 & n2491) | (n678 & n2492) | (n2491 & n2492);
  assign n2494 = n2490 | n2493;
  assign n2495 = x134 & ~n2494;
  assign n2496 = n937 & ~n963;
  assign n2497 = (~x132 & x133) | (~x132 & n880) | (x133 & n880);
  assign n2498 = (x132 & x133) | (x132 & n868) | (x133 & n868);
  assign n2499 = n2496 | n2498;
  assign n2500 = (n2496 & n2497) | (n2496 & n2499) | (n2497 & n2499);
  assign n2501 = x134 & ~n2500;
  assign n2502 = (~n2495 & n2500) | (~n2495 & n2501) | (n2500 & n2501);
  assign n2503 = x133 | n1231;
  assign n2504 = x133 & ~n2237;
  assign n2505 = (n678 & n2503) | (n678 & n2504) | (n2503 & n2504);
  assign n2506 = x133 | n1187;
  assign n2507 = (x132 & ~n763) | (x132 & n1097) | (~n763 & n1097);
  assign n2508 = x133 & n2507;
  assign n2509 = (~n763 & n2506) | (~n763 & n2508) | (n2506 & n2508);
  assign n2510 = n2505 | n2509;
  assign n2511 = ~n2226 & n2234;
  assign n2512 = (x132 & x133) | (x132 & n1012) | (x133 & n1012);
  assign n2513 = (x132 & ~x133) | (x132 & n1265) | (~x133 & n1265);
  assign n2514 = n2511 | n2513;
  assign n2515 = (n2511 & n2512) | (n2511 & n2514) | (n2512 & n2514);
  assign n2516 = x134 & ~n2515;
  assign n2517 = x134 & ~n2510;
  assign n2518 = (n2510 & ~n2516) | (n2510 & n2517) | (~n2516 & n2517);
  assign n2519 = (~x132 & x133) | (~x132 & n1323) | (x133 & n1323);
  assign n2520 = n2251 & n2519;
  assign n2521 = (x132 & ~x133) | (x132 & n1359) | (~x133 & n1359);
  assign n2522 = (x132 & x133) | (x132 & ~n1367) | (x133 & ~n1367);
  assign n2523 = ~n2520 & n2522;
  assign n2524 = (n2520 & n2521) | (n2520 & ~n2523) | (n2521 & ~n2523);
  assign n2525 = x134 & ~n2524;
  assign n2526 = (x132 & x133) | (x132 & ~n1340) | (x133 & ~n1340);
  assign n2527 = n2250 & ~n2526;
  assign n2528 = (~x132 & x133) | (~x132 & n1376) | (x133 & n1376);
  assign n2529 = (x132 & x133) | (x132 & n1384) | (x133 & n1384);
  assign n2530 = n2527 | n2529;
  assign n2531 = (n2527 & n2528) | (n2527 & n2530) | (n2528 & n2530);
  assign n2532 = x134 & ~n2531;
  assign n2533 = (~n2525 & n2531) | (~n2525 & n2532) | (n2531 & n2532);
  assign n2534 = (~x132 & x133) | (~x132 & n1396) | (x133 & n1396);
  assign n2535 = n2266 & n2534;
  assign n2536 = (x132 & ~x133) | (x132 & n1432) | (~x133 & n1432);
  assign n2537 = (x132 & x133) | (x132 & ~n1440) | (x133 & ~n1440);
  assign n2538 = ~n2535 & n2537;
  assign n2539 = (n2535 & n2536) | (n2535 & ~n2538) | (n2536 & ~n2538);
  assign n2540 = x134 & ~n2539;
  assign n2541 = (x132 & x133) | (x132 & ~n1413) | (x133 & ~n1413);
  assign n2542 = n2265 & ~n2541;
  assign n2543 = (~x132 & x133) | (~x132 & n1449) | (x133 & n1449);
  assign n2544 = (x132 & x133) | (x132 & n1457) | (x133 & n1457);
  assign n2545 = n2542 | n2544;
  assign n2546 = (n2542 & n2543) | (n2542 & n2545) | (n2543 & n2545);
  assign n2547 = x134 & ~n2546;
  assign n2548 = (~n2540 & n2546) | (~n2540 & n2547) | (n2546 & n2547);
  assign n2549 = (~x132 & x133) | (~x132 & n1469) | (x133 & n1469);
  assign n2550 = n2281 & n2549;
  assign n2551 = (x132 & ~x133) | (x132 & n1505) | (~x133 & n1505);
  assign n2552 = (x132 & x133) | (x132 & ~n1513) | (x133 & ~n1513);
  assign n2553 = ~n2550 & n2552;
  assign n2554 = (n2550 & n2551) | (n2550 & ~n2553) | (n2551 & ~n2553);
  assign n2555 = x134 & ~n2554;
  assign n2556 = (x132 & x133) | (x132 & ~n1486) | (x133 & ~n1486);
  assign n2557 = n2280 & ~n2556;
  assign n2558 = (~x132 & x133) | (~x132 & n1522) | (x133 & n1522);
  assign n2559 = (x132 & x133) | (x132 & n1530) | (x133 & n1530);
  assign n2560 = n2557 | n2559;
  assign n2561 = (n2557 & n2558) | (n2557 & n2560) | (n2558 & n2560);
  assign n2562 = x134 & ~n2561;
  assign n2563 = (~n2555 & n2561) | (~n2555 & n2562) | (n2561 & n2562);
  assign n2564 = (x132 & x133) | (x132 & n1558) | (x133 & n1558);
  assign n2565 = (~x132 & x133) | (~x132 & n1570) | (x133 & n1570);
  assign n2566 = n2564 & n2565;
  assign n2567 = (x132 & x133) | (x132 & ~n1598) | (x133 & ~n1598);
  assign n2568 = (x132 & ~x133) | (x132 & n1606) | (~x133 & n1606);
  assign n2569 = n2566 | n2568;
  assign n2570 = (n2566 & ~n2567) | (n2566 & n2569) | (~n2567 & n2569);
  assign n2571 = x134 & ~n2570;
  assign n2572 = (x132 & x133) | (x132 & ~n1550) | (x133 & ~n1550);
  assign n2573 = n2296 & ~n2572;
  assign n2574 = (~x132 & x133) | (~x132 & n1581) | (x133 & n1581);
  assign n2575 = (x132 & x133) | (x132 & n1589) | (x133 & n1589);
  assign n2576 = n2573 | n2575;
  assign n2577 = (n2573 & n2574) | (n2573 & n2576) | (n2574 & n2576);
  assign n2578 = x134 & ~n2577;
  assign n2579 = (~n2571 & n2577) | (~n2571 & n2578) | (n2577 & n2578);
  assign n2580 = (x132 & x133) | (x132 & n1635) | (x133 & n1635);
  assign n2581 = (~x132 & x133) | (~x132 & n1643) | (x133 & n1643);
  assign n2582 = n2580 & n2581;
  assign n2583 = (x132 & x133) | (x132 & ~n1671) | (x133 & ~n1671);
  assign n2584 = (x132 & ~x133) | (x132 & n1679) | (~x133 & n1679);
  assign n2585 = n2582 | n2584;
  assign n2586 = (n2582 & ~n2583) | (n2582 & n2585) | (~n2583 & n2585);
  assign n2587 = x134 & ~n2586;
  assign n2588 = (x132 & x133) | (x132 & ~n1626) | (x133 & ~n1626);
  assign n2589 = n2317 & ~n2588;
  assign n2590 = (~x132 & x133) | (~x132 & n1654) | (x133 & n1654);
  assign n2591 = (x132 & x133) | (x132 & n1662) | (x133 & n1662);
  assign n2592 = n2589 | n2591;
  assign n2593 = (n2589 & n2590) | (n2589 & n2592) | (n2590 & n2592);
  assign n2594 = x134 & ~n2593;
  assign n2595 = (~n2587 & n2593) | (~n2587 & n2594) | (n2593 & n2594);
  assign n2596 = (x132 & x133) | (x132 & n1708) | (x133 & n1708);
  assign n2597 = (~x132 & x133) | (~x132 & n1716) | (x133 & n1716);
  assign n2598 = n2596 & n2597;
  assign n2599 = (x132 & x133) | (x132 & ~n1744) | (x133 & ~n1744);
  assign n2600 = (x132 & ~x133) | (x132 & n1752) | (~x133 & n1752);
  assign n2601 = n2598 | n2600;
  assign n2602 = (n2598 & ~n2599) | (n2598 & n2601) | (~n2599 & n2601);
  assign n2603 = x134 & ~n2602;
  assign n2604 = (x132 & x133) | (x132 & ~n1699) | (x133 & ~n1699);
  assign n2605 = n2337 & ~n2604;
  assign n2606 = (~x132 & x133) | (~x132 & n1727) | (x133 & n1727);
  assign n2607 = (x132 & x133) | (x132 & n1735) | (x133 & n1735);
  assign n2608 = n2605 | n2607;
  assign n2609 = (n2605 & n2606) | (n2605 & n2608) | (n2606 & n2608);
  assign n2610 = x134 & ~n2609;
  assign n2611 = (~n2603 & n2609) | (~n2603 & n2610) | (n2609 & n2610);
  assign n2612 = (x132 & x133) | (x132 & n1807) | (x133 & n1807);
  assign n2613 = (~x132 & x133) | (~x132 & n1799) | (x133 & n1799);
  assign n2614 = n2612 & ~n2613;
  assign n2615 = x132 & n1789;
  assign n2616 = ~x132 & n1781;
  assign n2617 = (~x133 & n2615) | (~x133 & n2616) | (n2615 & n2616);
  assign n2618 = (n2612 & ~n2614) | (n2612 & n2617) | (~n2614 & n2617);
  assign n2619 = x134 & ~n2618;
  assign n2620 = (x132 & x133) | (x132 & ~n1816) | (x133 & ~n1816);
  assign n2621 = n2355 & ~n2620;
  assign n2622 = x133 | n2621;
  assign n2623 = (x132 & ~x133) | (x132 & n1772) | (~x133 & n1772);
  assign n2624 = (~x132 & n1764) | (~x132 & n2623) | (n1764 & n2623);
  assign n2625 = (n2621 & n2622) | (n2621 & n2623) | (n2622 & n2623);
  assign n2626 = (n2622 & n2624) | (n2622 & n2625) | (n2624 & n2625);
  assign n2627 = x134 & ~n2626;
  assign n2628 = (~n2619 & n2626) | (~n2619 & n2627) | (n2626 & n2627);
  assign n2629 = (x132 & x133) | (x132 & n1878) | (x133 & n1878);
  assign n2630 = (~x132 & x133) | (~x132 & n1870) | (x133 & n1870);
  assign n2631 = n2629 & ~n2630;
  assign n2632 = x132 & n1862;
  assign n2633 = ~x132 & n1854;
  assign n2634 = (~x133 & n2632) | (~x133 & n2633) | (n2632 & n2633);
  assign n2635 = (n2629 & ~n2631) | (n2629 & n2634) | (~n2631 & n2634);
  assign n2636 = x134 & ~n2635;
  assign n2637 = (x132 & x133) | (x132 & ~n1887) | (x133 & ~n1887);
  assign n2638 = n2373 & ~n2637;
  assign n2639 = x133 | n2638;
  assign n2640 = (x132 & ~x133) | (x132 & n1845) | (~x133 & n1845);
  assign n2641 = (~x132 & n1837) | (~x132 & n2640) | (n1837 & n2640);
  assign n2642 = (n2638 & n2639) | (n2638 & n2640) | (n2639 & n2640);
  assign n2643 = (n2639 & n2641) | (n2639 & n2642) | (n2641 & n2642);
  assign n2644 = x134 & ~n2643;
  assign n2645 = (~n2636 & n2643) | (~n2636 & n2644) | (n2643 & n2644);
  assign n2646 = (x132 & x133) | (x132 & n1946) | (x133 & n1946);
  assign n2647 = (~x132 & x133) | (~x132 & n1938) | (x133 & n1938);
  assign n2648 = n2646 & ~n2647;
  assign n2649 = x132 & n1915;
  assign n2650 = ~x132 & n1907;
  assign n2651 = (~x133 & n2649) | (~x133 & n2650) | (n2649 & n2650);
  assign n2652 = (n2646 & ~n2648) | (n2646 & n2651) | (~n2648 & n2651);
  assign n2653 = x134 & ~n2652;
  assign n2654 = (x132 & x133) | (x132 & ~n1955) | (x133 & ~n1955);
  assign n2655 = n2391 & ~n2654;
  assign n2656 = x133 | n2655;
  assign n2657 = (x132 & ~x133) | (x132 & n1924) | (~x133 & n1924);
  assign n2658 = (~x132 & n1930) | (~x132 & n2657) | (n1930 & n2657);
  assign n2659 = (n2655 & n2656) | (n2655 & n2657) | (n2656 & n2657);
  assign n2660 = (n2656 & n2658) | (n2656 & n2659) | (n2658 & n2659);
  assign n2661 = x134 & ~n2660;
  assign n2662 = (~n2653 & n2660) | (~n2653 & n2661) | (n2660 & n2661);
  assign n2663 = (x132 & x133) | (x132 & n2015) | (x133 & n2015);
  assign n2664 = (~x132 & x133) | (~x132 & n2007) | (x133 & n2007);
  assign n2665 = n2663 & ~n2664;
  assign n2666 = x132 & n1984;
  assign n2667 = ~x132 & n1976;
  assign n2668 = (~x133 & n2666) | (~x133 & n2667) | (n2666 & n2667);
  assign n2669 = (n2663 & ~n2665) | (n2663 & n2668) | (~n2665 & n2668);
  assign n2670 = x134 & ~n2669;
  assign n2671 = (x132 & x133) | (x132 & ~n2024) | (x133 & ~n2024);
  assign n2672 = n2409 & ~n2671;
  assign n2673 = x133 | n2672;
  assign n2674 = (x132 & ~x133) | (x132 & n1993) | (~x133 & n1993);
  assign n2675 = (~x132 & n1999) | (~x132 & n2674) | (n1999 & n2674);
  assign n2676 = (n2672 & n2673) | (n2672 & n2674) | (n2673 & n2674);
  assign n2677 = (n2673 & n2675) | (n2673 & n2676) | (n2675 & n2676);
  assign n2678 = x134 & ~n2677;
  assign n2679 = (~n2670 & n2677) | (~n2670 & n2678) | (n2677 & n2678);
  assign n2680 = (x132 & x133) | (x132 & n2084) | (x133 & n2084);
  assign n2681 = (~x132 & x133) | (~x132 & n2076) | (x133 & n2076);
  assign n2682 = n2680 & ~n2681;
  assign n2683 = x132 & n2053;
  assign n2684 = ~x132 & n2045;
  assign n2685 = (~x133 & n2683) | (~x133 & n2684) | (n2683 & n2684);
  assign n2686 = (n2680 & ~n2682) | (n2680 & n2685) | (~n2682 & n2685);
  assign n2687 = x134 & ~n2686;
  assign n2688 = (x132 & x133) | (x132 & ~n2093) | (x133 & ~n2093);
  assign n2689 = n2427 & ~n2688;
  assign n2690 = x133 | n2689;
  assign n2691 = (x132 & ~x133) | (x132 & n2062) | (~x133 & n2062);
  assign n2692 = (~x132 & n2068) | (~x132 & n2691) | (n2068 & n2691);
  assign n2693 = (n2689 & n2690) | (n2689 & n2691) | (n2690 & n2691);
  assign n2694 = (n2690 & n2692) | (n2690 & n2693) | (n2692 & n2693);
  assign n2695 = x134 & ~n2694;
  assign n2696 = (~n2687 & n2694) | (~n2687 & n2695) | (n2694 & n2695);
  assign n2697 = (x132 & x133) | (x132 & ~n2120) | (x133 & ~n2120);
  assign n2698 = (x132 & ~x133) | (x132 & n2114) | (~x133 & n2114);
  assign n2699 = ~n2697 & n2698;
  assign n2700 = (x132 & x133) | (x132 & n2152) | (x133 & n2152);
  assign n2701 = (~x132 & x133) | (~x132 & n2144) | (x133 & n2144);
  assign n2702 = n2700 & ~n2701;
  assign n2703 = (n2699 & n2700) | (n2699 & ~n2702) | (n2700 & ~n2702);
  assign n2704 = x134 & ~n2703;
  assign n2705 = (x132 & x133) | (x132 & ~n2161) | (x133 & ~n2161);
  assign n2706 = n2444 & ~n2705;
  assign n2707 = x133 | n2706;
  assign n2708 = (x132 & ~x133) | (x132 & n2129) | (~x133 & n2129);
  assign n2709 = (~x132 & n2135) | (~x132 & n2708) | (n2135 & n2708);
  assign n2710 = (n2706 & n2707) | (n2706 & n2708) | (n2707 & n2708);
  assign n2711 = (n2707 & n2709) | (n2707 & n2710) | (n2709 & n2710);
  assign n2712 = x134 & ~n2711;
  assign n2713 = (~n2704 & n2711) | (~n2704 & n2712) | (n2711 & n2712);
  assign n2714 = x133 | n222;
  assign n2715 = x133 & n404;
  assign n2716 = (~n763 & n2714) | (~n763 & n2715) | (n2714 & n2715);
  assign n2717 = x133 | n267;
  assign n2718 = x133 & ~n2455;
  assign n2719 = (n678 & n2717) | (n678 & n2718) | (n2717 & n2718);
  assign n2720 = n2716 | n2719;
  assign n2721 = x134 & ~n2720;
  assign n2722 = n2174 & ~n2178;
  assign n2723 = (~x132 & x133) | (~x132 & n178) | (x133 & n178);
  assign n2724 = (x132 & x133) | (x132 & n492) | (x133 & n492);
  assign n2725 = n2722 | n2724;
  assign n2726 = (n2722 & n2723) | (n2722 & n2725) | (n2723 & n2725);
  assign n2727 = x134 & ~n2726;
  assign n2728 = (~n2721 & n2726) | (~n2721 & n2727) | (n2726 & n2727);
  assign n2729 = (x132 & x133) | (x132 & n674) | (x133 & n674);
  assign n2730 = (~x132 & x133) | (~x132 & n806) | (x133 & n806);
  assign n2731 = n2729 & ~n2730;
  assign n2732 = x132 & n630;
  assign n2733 = ~x132 & n585;
  assign n2734 = (~x133 & n2732) | (~x133 & n2733) | (n2732 & n2733);
  assign n2735 = (n2729 & ~n2731) | (n2729 & n2734) | (~n2731 & n2734);
  assign n2736 = x134 & ~n2735;
  assign n2737 = (x133 & n2201) | (x133 & n2202) | (n2201 & n2202);
  assign n2738 = (x132 & x133) | (x132 & ~n759) | (x133 & ~n759);
  assign n2739 = n2472 | n2737;
  assign n2740 = (n2737 & ~n2738) | (n2737 & n2739) | (~n2738 & n2739);
  assign n2741 = x134 & ~n2740;
  assign n2742 = (~n2736 & n2740) | (~n2736 & n2741) | (n2740 & n2741);
  assign n2743 = (x132 & x133) | (x132 & n905) | (x133 & n905);
  assign n2744 = (~x132 & x133) | (~x132 & n950) | (x133 & n950);
  assign n2745 = n2743 & ~n2744;
  assign n2746 = x132 & n893;
  assign n2747 = ~x132 & n880;
  assign n2748 = (~x133 & n2746) | (~x133 & n2747) | (n2746 & n2747);
  assign n2749 = (n2743 & ~n2745) | (n2743 & n2748) | (~n2745 & n2748);
  assign n2750 = x134 & ~n2749;
  assign n2751 = (x133 & n2218) | (x133 & n2219) | (n2218 & n2219);
  assign n2752 = (x132 & x133) | (x132 & ~n936) | (x133 & ~n936);
  assign n2753 = n2488 | n2751;
  assign n2754 = (n2751 & ~n2752) | (n2751 & n2753) | (~n2752 & n2753);
  assign n2755 = x134 & ~n2754;
  assign n2756 = (~n2750 & n2754) | (~n2750 & n2755) | (n2754 & n2755);
  assign n2757 = x133 | n1140;
  assign n2758 = n1012 & ~n1013;
  assign n2759 = (n678 & n2757) | (n678 & n2758) | (n2757 & n2758);
  assign n2760 = n1310 & n2226;
  assign n2761 = (~n763 & n1098) | (~n763 & n2760) | (n1098 & n2760);
  assign n2762 = n2759 | n2761;
  assign n2763 = x134 & ~n2762;
  assign n2764 = (x132 & x133) | (x132 & n1231) | (x133 & n1231);
  assign n2765 = (x132 & x133) | (x132 & ~n1187) | (x133 & ~n1187);
  assign n2766 = n2513 & ~n2765;
  assign n2767 = (~x132 & x133) | (~x132 & n1054) | (x133 & n1054);
  assign n2768 = n2764 & ~n2767;
  assign n2769 = (n2764 & n2766) | (n2764 & ~n2768) | (n2766 & ~n2768);
  assign n2770 = x134 & ~n2769;
  assign n2771 = (~n2763 & n2769) | (~n2763 & n2770) | (n2769 & n2770);
  assign n2772 = x133 | n1348;
  assign n2773 = x133 & ~n2526;
  assign n2774 = (n678 & n2772) | (n678 & n2773) | (n2772 & n2773);
  assign n2775 = x133 | n1323;
  assign n2776 = x133 & n1385;
  assign n2777 = (~n763 & n2775) | (~n763 & n2776) | (n2775 & n2776);
  assign n2778 = n2774 | n2777;
  assign n2779 = x133 & n1332;
  assign n2780 = x133 | n1376;
  assign n2781 = (~n763 & n2779) | (~n763 & n2780) | (n2779 & n2780);
  assign n2782 = x133 | n1359;
  assign n2783 = x133 & ~n2522;
  assign n2784 = (n678 & n2782) | (n678 & n2783) | (n2782 & n2783);
  assign n2785 = n2781 | n2784;
  assign n2786 = x134 & ~n2785;
  assign n2787 = x134 & ~n2778;
  assign n2788 = (n2778 & ~n2786) | (n2778 & n2787) | (~n2786 & n2787);
  assign n2789 = x133 | n1421;
  assign n2790 = x133 & ~n2541;
  assign n2791 = (n678 & n2789) | (n678 & n2790) | (n2789 & n2790);
  assign n2792 = x133 | n1396;
  assign n2793 = (x132 & ~n763) | (x132 & n1457) | (~n763 & n1457);
  assign n2794 = x133 & n2793;
  assign n2795 = (~n763 & n2792) | (~n763 & n2794) | (n2792 & n2794);
  assign n2796 = n2791 | n2795;
  assign n2797 = x133 & n1405;
  assign n2798 = x133 | n1449;
  assign n2799 = (~n763 & n2797) | (~n763 & n2798) | (n2797 & n2798);
  assign n2800 = x133 | n1432;
  assign n2801 = x133 & ~n2537;
  assign n2802 = (n678 & n2800) | (n678 & n2801) | (n2800 & n2801);
  assign n2803 = n2799 | n2802;
  assign n2804 = x134 & ~n2803;
  assign n2805 = x134 & ~n2796;
  assign n2806 = (n2796 & ~n2804) | (n2796 & n2805) | (~n2804 & n2805);
  assign n2807 = x133 | n1494;
  assign n2808 = x133 & ~n2556;
  assign n2809 = (n678 & n2807) | (n678 & n2808) | (n2807 & n2808);
  assign n2810 = x133 | n1469;
  assign n2811 = (x132 & ~n763) | (x132 & n1530) | (~n763 & n1530);
  assign n2812 = x133 & n2811;
  assign n2813 = (~n763 & n2810) | (~n763 & n2812) | (n2810 & n2812);
  assign n2814 = n2809 | n2813;
  assign n2815 = x133 & n1478;
  assign n2816 = x133 | n1522;
  assign n2817 = (~n763 & n2815) | (~n763 & n2816) | (n2815 & n2816);
  assign n2818 = x133 | n1505;
  assign n2819 = x133 & ~n2552;
  assign n2820 = (n678 & n2818) | (n678 & n2819) | (n2818 & n2819);
  assign n2821 = n2817 | n2820;
  assign n2822 = x134 & ~n2821;
  assign n2823 = x134 & ~n2814;
  assign n2824 = (n2814 & ~n2822) | (n2814 & n2823) | (~n2822 & n2823);
  assign n2825 = n2288 & ~n2292;
  assign n2826 = (~x132 & x133) | (~x132 & n1558) | (x133 & n1558);
  assign n2827 = (x132 & x133) | (x132 & n1598) | (x133 & n1598);
  assign n2828 = n2825 | n2827;
  assign n2829 = (n2825 & n2826) | (n2825 & n2828) | (n2826 & n2828);
  assign n2830 = x134 & ~n2829;
  assign n2831 = n1543 & n1590;
  assign n2832 = (n2565 & ~n2572) | (n2565 & n2831) | (~n2572 & n2831);
  assign n2833 = n2831 | n2832;
  assign n2834 = x134 & ~n2833;
  assign n2835 = (~n2830 & n2833) | (~n2830 & n2834) | (n2833 & n2834);
  assign n2836 = n2308 & ~n2312;
  assign n2837 = (~x132 & x133) | (~x132 & n1635) | (x133 & n1635);
  assign n2838 = (x132 & x133) | (x132 & n1671) | (x133 & n1671);
  assign n2839 = n2836 | n2838;
  assign n2840 = (n2836 & n2837) | (n2836 & n2839) | (n2837 & n2839);
  assign n2841 = x134 & ~n2840;
  assign n2842 = n1619 & n1663;
  assign n2843 = (n2581 & ~n2588) | (n2581 & n2842) | (~n2588 & n2842);
  assign n2844 = n2842 | n2843;
  assign n2845 = x134 & ~n2844;
  assign n2846 = (~n2841 & n2844) | (~n2841 & n2845) | (n2844 & n2845);
  assign n2847 = n2328 & ~n2332;
  assign n2848 = (~x132 & x133) | (~x132 & n1708) | (x133 & n1708);
  assign n2849 = (x132 & x133) | (x132 & n1744) | (x133 & n1744);
  assign n2850 = n2847 | n2849;
  assign n2851 = (n2847 & n2848) | (n2847 & n2850) | (n2848 & n2850);
  assign n2852 = x134 & ~n2851;
  assign n2853 = n1692 & n1736;
  assign n2854 = (n2597 & ~n2604) | (n2597 & n2853) | (~n2604 & n2853);
  assign n2855 = n2853 | n2854;
  assign n2856 = x134 & ~n2855;
  assign n2857 = (~n2852 & n2855) | (~n2852 & n2856) | (n2855 & n2856);
  assign n2858 = x133 | n1824;
  assign n2859 = x133 & ~n2620;
  assign n2860 = (n678 & n2858) | (n678 & n2859) | (n2858 & n2859);
  assign n2861 = x133 | n1799;
  assign n2862 = (x132 & ~n763) | (x132 & n1764) | (~n763 & n1764);
  assign n2863 = x133 & n2862;
  assign n2864 = (~n763 & n2861) | (~n763 & n2863) | (n2861 & n2863);
  assign n2865 = n2860 | n2864;
  assign n2866 = (x132 & x133) | (x132 & ~n1781) | (x133 & ~n1781);
  assign n2867 = n2623 & ~n2866;
  assign n2868 = (~x132 & x133) | (~x132 & n1807) | (x133 & n1807);
  assign n2869 = (x132 & x133) | (x132 & n1789) | (x133 & n1789);
  assign n2870 = n2868 & ~n2869;
  assign n2871 = (n2867 & n2868) | (n2867 & ~n2870) | (n2868 & ~n2870);
  assign n2872 = x134 & ~n2871;
  assign n2873 = x134 & ~n2865;
  assign n2874 = (n2865 & ~n2872) | (n2865 & n2873) | (~n2872 & n2873);
  assign n2875 = x133 | n1894;
  assign n2876 = x133 & ~n2637;
  assign n2877 = (n678 & n2875) | (n678 & n2876) | (n2875 & n2876);
  assign n2878 = x133 | n1870;
  assign n2879 = (x132 & ~n763) | (x132 & n1837) | (~n763 & n1837);
  assign n2880 = x133 & n2879;
  assign n2881 = (~n763 & n2878) | (~n763 & n2880) | (n2878 & n2880);
  assign n2882 = n2877 | n2881;
  assign n2883 = (x132 & x133) | (x132 & ~n1854) | (x133 & ~n1854);
  assign n2884 = n2640 & ~n2883;
  assign n2885 = (~x132 & x133) | (~x132 & n1878) | (x133 & n1878);
  assign n2886 = (x132 & x133) | (x132 & n1862) | (x133 & n1862);
  assign n2887 = n2885 & ~n2886;
  assign n2888 = (n2884 & n2885) | (n2884 & ~n2887) | (n2885 & ~n2887);
  assign n2889 = x134 & ~n2888;
  assign n2890 = x134 & ~n2882;
  assign n2891 = (n2882 & ~n2889) | (n2882 & n2890) | (~n2889 & n2890);
  assign n2892 = x133 | n1963;
  assign n2893 = x133 & ~n2654;
  assign n2894 = (n678 & n2892) | (n678 & n2893) | (n2892 & n2893);
  assign n2895 = x133 | n1938;
  assign n2896 = (x132 & ~n763) | (x132 & n1930) | (~n763 & n1930);
  assign n2897 = x133 & n2896;
  assign n2898 = (~n763 & n2895) | (~n763 & n2897) | (n2895 & n2897);
  assign n2899 = n2894 | n2898;
  assign n2900 = (x132 & x133) | (x132 & ~n1907) | (x133 & ~n1907);
  assign n2901 = n2657 & ~n2900;
  assign n2902 = (~x132 & x133) | (~x132 & n1946) | (x133 & n1946);
  assign n2903 = (x132 & x133) | (x132 & n1915) | (x133 & n1915);
  assign n2904 = n2902 & ~n2903;
  assign n2905 = (n2901 & n2902) | (n2901 & ~n2904) | (n2902 & ~n2904);
  assign n2906 = x134 & ~n2905;
  assign n2907 = x134 & ~n2899;
  assign n2908 = (n2899 & ~n2906) | (n2899 & n2907) | (~n2906 & n2907);
  assign n2909 = x133 | n2032;
  assign n2910 = x133 & ~n2671;
  assign n2911 = (n678 & n2909) | (n678 & n2910) | (n2909 & n2910);
  assign n2912 = x133 | n2007;
  assign n2913 = (x132 & ~n763) | (x132 & n1999) | (~n763 & n1999);
  assign n2914 = x133 & n2913;
  assign n2915 = (~n763 & n2912) | (~n763 & n2914) | (n2912 & n2914);
  assign n2916 = n2911 | n2915;
  assign n2917 = (x132 & x133) | (x132 & ~n1976) | (x133 & ~n1976);
  assign n2918 = n2674 & ~n2917;
  assign n2919 = (~x132 & x133) | (~x132 & n2015) | (x133 & n2015);
  assign n2920 = (x132 & x133) | (x132 & n1984) | (x133 & n1984);
  assign n2921 = n2919 & ~n2920;
  assign n2922 = (n2918 & n2919) | (n2918 & ~n2921) | (n2919 & ~n2921);
  assign n2923 = x134 & ~n2922;
  assign n2924 = x134 & ~n2916;
  assign n2925 = (n2916 & ~n2923) | (n2916 & n2924) | (~n2923 & n2924);
  assign n2926 = x133 | n2101;
  assign n2927 = x133 & ~n2688;
  assign n2928 = (n678 & n2926) | (n678 & n2927) | (n2926 & n2927);
  assign n2929 = x133 | n2076;
  assign n2930 = (x132 & ~n763) | (x132 & n2068) | (~n763 & n2068);
  assign n2931 = x133 & n2930;
  assign n2932 = (~n763 & n2929) | (~n763 & n2931) | (n2929 & n2931);
  assign n2933 = n2928 | n2932;
  assign n2934 = (x132 & x133) | (x132 & ~n2045) | (x133 & ~n2045);
  assign n2935 = n2691 & ~n2934;
  assign n2936 = (~x132 & x133) | (~x132 & n2084) | (x133 & n2084);
  assign n2937 = (x132 & x133) | (x132 & n2053) | (x133 & n2053);
  assign n2938 = n2936 & ~n2937;
  assign n2939 = (n2935 & n2936) | (n2935 & ~n2938) | (n2936 & ~n2938);
  assign n2940 = x134 & ~n2939;
  assign n2941 = x134 & ~n2933;
  assign n2942 = (n2933 & ~n2940) | (n2933 & n2941) | (~n2940 & n2941);
  assign n2943 = x133 | n2166;
  assign n2944 = x133 & ~n2705;
  assign n2945 = (n678 & n2943) | (n678 & n2944) | (n2943 & n2944);
  assign n2946 = x133 | n2144;
  assign n2947 = (x132 & ~n763) | (x132 & n2135) | (~n763 & n2135);
  assign n2948 = x133 & n2947;
  assign n2949 = (~n763 & n2946) | (~n763 & n2948) | (n2946 & n2948);
  assign n2950 = n2945 | n2949;
  assign n2951 = (x132 & x133) | (x132 & ~n2114) | (x133 & ~n2114);
  assign n2952 = n2708 & ~n2951;
  assign n2953 = x133 | n2952;
  assign n2954 = (~x132 & n2120) | (~x132 & n2153) | (n2120 & n2153);
  assign n2955 = (n2153 & n2952) | (n2153 & n2953) | (n2952 & n2953);
  assign n2956 = (n2953 & n2954) | (n2953 & n2955) | (n2954 & n2955);
  assign n2957 = x134 & ~n2956;
  assign n2958 = x134 & ~n2950;
  assign n2959 = (n2950 & ~n2957) | (n2950 & n2958) | (~n2957 & n2958);
  assign n2960 = (n496 & n497) | (n496 & ~n498) | (n497 & ~n498);
  assign n2961 = (n854 & n855) | (n854 & ~n856) | (n855 & ~n856);
  assign n2962 = (n966 & n967) | (n966 & ~n968) | (n967 & ~n968);
  assign n2963 = (n1313 & n1314) | (n1313 & ~n1315) | (n1314 & ~n1315);
  assign n2964 = (n1351 & n1352) | (n1351 & ~n1388) | (n1352 & ~n1388);
  assign n2965 = (n1424 & n1425) | (n1424 & ~n1461) | (n1425 & ~n1461);
  assign n2966 = (n1497 & n1498) | (n1497 & ~n1534) | (n1498 & ~n1534);
  assign n2967 = (n1573 & n1574) | (n1573 & ~n1610) | (n1574 & ~n1610);
  assign n2968 = (n1646 & n1647) | (n1646 & ~n1683) | (n1647 & ~n1683);
  assign n2969 = (n1719 & n1720) | (n1719 & ~n1756) | (n1720 & ~n1756);
  assign n2970 = (n1827 & n1828) | (n1827 & ~n1829) | (n1828 & ~n1829);
  assign n2971 = (n1897 & n1898) | (n1897 & ~n1899) | (n1898 & ~n1899);
  assign n2972 = (n1966 & n1967) | (n1966 & ~n1968) | (n1967 & ~n1968);
  assign n2973 = (n2035 & n2036) | (n2035 & ~n2037) | (n2036 & ~n2037);
  assign n2974 = (n2104 & n2105) | (n2104 & ~n2106) | (n2105 & ~n2106);
  assign n2975 = (n2169 & n2170) | (n2169 & ~n2171) | (n2170 & ~n2171);
  assign n2976 = (n2181 & n2182) | (n2181 & ~n2190) | (n2182 & ~n2190);
  assign n2977 = (n2198 & n2199) | (n2198 & ~n2207) | (n2199 & ~n2207);
  assign n2978 = (n2215 & n2216) | (n2215 & ~n2224) | (n2216 & ~n2224);
  assign n2979 = (n2231 & n2232) | (n2231 & ~n2240) | (n2232 & ~n2240);
  assign n2980 = (n2253 & n2254) | (n2253 & ~n2255) | (n2254 & ~n2255);
  assign n2981 = (n2268 & n2269) | (n2268 & ~n2270) | (n2269 & ~n2270);
  assign n2982 = (n2283 & n2284) | (n2283 & ~n2285) | (n2284 & ~n2285);
  assign n2983 = (n2303 & n2304) | (n2303 & ~n2305) | (n2304 & ~n2305);
  assign n2984 = (n2323 & n2324) | (n2323 & ~n2325) | (n2324 & ~n2325);
  assign n2985 = (n2343 & n2344) | (n2343 & ~n2345) | (n2344 & ~n2345);
  assign n2986 = (n2361 & n2362) | (n2361 & ~n2363) | (n2362 & ~n2363);
  assign n2987 = (n2379 & n2380) | (n2379 & ~n2381) | (n2380 & ~n2381);
  assign n2988 = (n2397 & n2398) | (n2397 & ~n2399) | (n2398 & ~n2399);
  assign n2989 = (n2415 & n2416) | (n2415 & ~n2417) | (n2416 & ~n2417);
  assign n2990 = (n2433 & n2434) | (n2433 & ~n2435) | (n2434 & ~n2435);
  assign n2991 = (n2451 & n2452) | (n2451 & ~n2453) | (n2452 & ~n2453);
  assign n2992 = (n2460 & n2461) | (n2460 & ~n2469) | (n2461 & ~n2469);
  assign n2993 = (n2478 & n2479) | (n2478 & ~n2485) | (n2479 & ~n2485);
  assign n2994 = (n2494 & n2495) | (n2494 & ~n2501) | (n2495 & ~n2501);
  assign n2995 = (n2515 & n2516) | (n2515 & ~n2517) | (n2516 & ~n2517);
  assign n2996 = (n2524 & n2525) | (n2524 & ~n2532) | (n2525 & ~n2532);
  assign n2997 = (n2539 & n2540) | (n2539 & ~n2547) | (n2540 & ~n2547);
  assign n2998 = (n2554 & n2555) | (n2554 & ~n2562) | (n2555 & ~n2562);
  assign n2999 = (n2570 & n2571) | (n2570 & ~n2578) | (n2571 & ~n2578);
  assign n3000 = (n2586 & n2587) | (n2586 & ~n2594) | (n2587 & ~n2594);
  assign n3001 = (n2602 & n2603) | (n2602 & ~n2610) | (n2603 & ~n2610);
  assign n3002 = (n2618 & n2619) | (n2618 & ~n2627) | (n2619 & ~n2627);
  assign n3003 = (n2635 & n2636) | (n2635 & ~n2644) | (n2636 & ~n2644);
  assign n3004 = (n2652 & n2653) | (n2652 & ~n2661) | (n2653 & ~n2661);
  assign n3005 = (n2669 & n2670) | (n2669 & ~n2678) | (n2670 & ~n2678);
  assign n3006 = (n2686 & n2687) | (n2686 & ~n2695) | (n2687 & ~n2695);
  assign n3007 = (n2703 & n2704) | (n2703 & ~n2712) | (n2704 & ~n2712);
  assign n3008 = (n2720 & n2721) | (n2720 & ~n2727) | (n2721 & ~n2727);
  assign n3009 = (n2735 & n2736) | (n2735 & ~n2741) | (n2736 & ~n2741);
  assign n3010 = (n2749 & n2750) | (n2749 & ~n2755) | (n2750 & ~n2755);
  assign n3011 = (n2762 & n2763) | (n2762 & ~n2770) | (n2763 & ~n2770);
  assign n3012 = (n2785 & n2786) | (n2785 & ~n2787) | (n2786 & ~n2787);
  assign n3013 = (n2803 & n2804) | (n2803 & ~n2805) | (n2804 & ~n2805);
  assign n3014 = (n2821 & n2822) | (n2821 & ~n2823) | (n2822 & ~n2823);
  assign n3015 = (n2829 & n2830) | (n2829 & ~n2834) | (n2830 & ~n2834);
  assign n3016 = (n2840 & n2841) | (n2840 & ~n2845) | (n2841 & ~n2845);
  assign n3017 = (n2851 & n2852) | (n2851 & ~n2856) | (n2852 & ~n2856);
  assign n3018 = (n2871 & n2872) | (n2871 & ~n2873) | (n2872 & ~n2873);
  assign n3019 = (n2888 & n2889) | (n2888 & ~n2890) | (n2889 & ~n2890);
  assign n3020 = (n2905 & n2906) | (n2905 & ~n2907) | (n2906 & ~n2907);
  assign n3021 = (n2922 & n2923) | (n2922 & ~n2924) | (n2923 & ~n2924);
  assign n3022 = (n2939 & n2940) | (n2939 & ~n2941) | (n2940 & ~n2941);
  assign n3023 = (n2956 & n2957) | (n2956 & ~n2958) | (n2957 & ~n2958);
  assign y0 = n499;
  assign y1 = n857;
  assign y2 = n969;
  assign y3 = n1316;
  assign y4 = n1389;
  assign y5 = n1462;
  assign y6 = n1535;
  assign y7 = n1611;
  assign y8 = n1684;
  assign y9 = n1757;
  assign y10 = n1830;
  assign y11 = n1900;
  assign y12 = n1969;
  assign y13 = n2038;
  assign y14 = n2107;
  assign y15 = n2172;
  assign y16 = n2191;
  assign y17 = n2208;
  assign y18 = n2225;
  assign y19 = n2241;
  assign y20 = n2256;
  assign y21 = n2271;
  assign y22 = n2286;
  assign y23 = n2306;
  assign y24 = n2326;
  assign y25 = n2346;
  assign y26 = n2364;
  assign y27 = n2382;
  assign y28 = n2400;
  assign y29 = n2418;
  assign y30 = n2436;
  assign y31 = n2454;
  assign y32 = n2470;
  assign y33 = n2486;
  assign y34 = n2502;
  assign y35 = n2518;
  assign y36 = n2533;
  assign y37 = n2548;
  assign y38 = n2563;
  assign y39 = n2579;
  assign y40 = n2595;
  assign y41 = n2611;
  assign y42 = n2628;
  assign y43 = n2645;
  assign y44 = n2662;
  assign y45 = n2679;
  assign y46 = n2696;
  assign y47 = n2713;
  assign y48 = n2728;
  assign y49 = n2742;
  assign y50 = n2756;
  assign y51 = n2771;
  assign y52 = n2788;
  assign y53 = n2806;
  assign y54 = n2824;
  assign y55 = n2835;
  assign y56 = n2846;
  assign y57 = n2857;
  assign y58 = n2874;
  assign y59 = n2891;
  assign y60 = n2908;
  assign y61 = n2925;
  assign y62 = n2942;
  assign y63 = n2959;
  assign y64 = n2960;
  assign y65 = n2961;
  assign y66 = n2962;
  assign y67 = n2963;
  assign y68 = n2964;
  assign y69 = n2965;
  assign y70 = n2966;
  assign y71 = n2967;
  assign y72 = n2968;
  assign y73 = n2969;
  assign y74 = n2970;
  assign y75 = n2971;
  assign y76 = n2972;
  assign y77 = n2973;
  assign y78 = n2974;
  assign y79 = n2975;
  assign y80 = n2976;
  assign y81 = n2977;
  assign y82 = n2978;
  assign y83 = n2979;
  assign y84 = n2980;
  assign y85 = n2981;
  assign y86 = n2982;
  assign y87 = n2983;
  assign y88 = n2984;
  assign y89 = n2985;
  assign y90 = n2986;
  assign y91 = n2987;
  assign y92 = n2988;
  assign y93 = n2989;
  assign y94 = n2990;
  assign y95 = n2991;
  assign y96 = n2992;
  assign y97 = n2993;
  assign y98 = n2994;
  assign y99 = n2995;
  assign y100 = n2996;
  assign y101 = n2997;
  assign y102 = n2998;
  assign y103 = n2999;
  assign y104 = n3000;
  assign y105 = n3001;
  assign y106 = n3002;
  assign y107 = n3003;
  assign y108 = n3004;
  assign y109 = n3005;
  assign y110 = n3006;
  assign y111 = n3007;
  assign y112 = n3008;
  assign y113 = n3009;
  assign y114 = n3010;
  assign y115 = n3011;
  assign y116 = n3012;
  assign y117 = n3013;
  assign y118 = n3014;
  assign y119 = n3015;
  assign y120 = n3016;
  assign y121 = n3017;
  assign y122 = n3018;
  assign y123 = n3019;
  assign y124 = n3020;
  assign y125 = n3021;
  assign y126 = n3022;
  assign y127 = n3023;
endmodule

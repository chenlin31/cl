// Benchmark "top" written by ABC on Wed Jun 26 20:37:56 2019

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] ,
    \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] ,
    \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] ,
    \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] ,
    \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] ,
    \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] ,
    \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] , \b[60] ,
    \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] , \b[68] ,
    \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] , \b[76] ,
    \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] , \b[84] ,
    \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] ,
    \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127] , cOut  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] ,
    \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] ,
    \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] ,
    \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] ,
    \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] ,
    \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] ,
    \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] ,
    \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] ,
    \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] ,
    \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] ,
    \b[76] , \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] ,
    \b[84] , \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] ,
    \b[92] , \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] , cOut;
  wire new_n386_, new_n387_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n431_, new_n432_, new_n433_, new_n434_,
    new_n435_, new_n436_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1012_, new_n1013_, new_n1014_, new_n1015_,
    new_n1016_, new_n1017_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1075_, new_n1076_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1089_, new_n1090_, new_n1091_, new_n1092_,
    new_n1093_, new_n1094_, new_n1096_, new_n1097_, new_n1098_, new_n1099_,
    new_n1100_, new_n1101_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1117_, new_n1118_, new_n1119_, new_n1120_,
    new_n1121_, new_n1122_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1138_, new_n1139_, new_n1140_, new_n1141_,
    new_n1142_, new_n1143_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1159_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1180_, new_n1181_, new_n1182_, new_n1183_,
    new_n1184_, new_n1185_, new_n1187_, new_n1188_, new_n1189_, new_n1190_,
    new_n1191_, new_n1192_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1222_, new_n1223_, new_n1224_, new_n1225_,
    new_n1226_, new_n1227_, new_n1229_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1234_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_, new_n1241_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1254_, new_n1255_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1264_, new_n1265_, new_n1266_, new_n1267_,
    new_n1268_, new_n1269_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_;
  assign new_n386_ = \a[0]  & \b[0] ;
  assign new_n387_ = ~\a[0]  & ~\b[0] ;
  assign \f[0]  = ~new_n386_ & ~new_n387_;
  assign new_n389_ = ~\a[1]  & ~\b[1] ;
  assign new_n390_ = \a[1]  & \b[1] ;
  assign new_n391_ = ~new_n389_ & ~new_n390_;
  assign new_n392_ = new_n386_ & ~new_n391_;
  assign new_n393_ = ~new_n386_ & new_n391_;
  assign \f[1]  = new_n392_ | new_n393_;
  assign new_n395_ = ~\a[2]  & ~\b[2] ;
  assign new_n396_ = \a[2]  & \b[2] ;
  assign new_n397_ = ~new_n395_ & ~new_n396_;
  assign new_n398_ = ~new_n386_ & ~new_n390_;
  assign new_n399_ = ~new_n389_ & ~new_n398_;
  assign new_n400_ = ~new_n397_ & ~new_n399_;
  assign new_n401_ = new_n397_ & new_n399_;
  assign \f[2]  = ~new_n400_ & ~new_n401_;
  assign new_n403_ = ~\a[3]  & ~\b[3] ;
  assign new_n404_ = \a[3]  & \b[3] ;
  assign new_n405_ = ~new_n403_ & ~new_n404_;
  assign new_n406_ = ~new_n396_ & ~new_n401_;
  assign new_n407_ = ~new_n405_ & new_n406_;
  assign new_n408_ = new_n405_ & ~new_n406_;
  assign \f[3]  = ~new_n407_ & ~new_n408_;
  assign new_n410_ = ~\a[4]  & ~\b[4] ;
  assign new_n411_ = \a[4]  & \b[4] ;
  assign new_n412_ = ~new_n410_ & ~new_n411_;
  assign new_n413_ = ~new_n404_ & ~new_n408_;
  assign new_n414_ = ~new_n412_ & new_n413_;
  assign new_n415_ = new_n412_ & ~new_n413_;
  assign \f[4]  = ~new_n414_ & ~new_n415_;
  assign new_n417_ = ~\a[5]  & ~\b[5] ;
  assign new_n418_ = \a[5]  & \b[5] ;
  assign new_n419_ = ~new_n417_ & ~new_n418_;
  assign new_n420_ = ~new_n411_ & ~new_n415_;
  assign new_n421_ = ~new_n419_ & new_n420_;
  assign new_n422_ = new_n419_ & ~new_n420_;
  assign \f[5]  = ~new_n421_ & ~new_n422_;
  assign new_n424_ = ~\a[6]  & ~\b[6] ;
  assign new_n425_ = \a[6]  & \b[6] ;
  assign new_n426_ = ~new_n424_ & ~new_n425_;
  assign new_n427_ = ~new_n418_ & ~new_n422_;
  assign new_n428_ = ~new_n426_ & new_n427_;
  assign new_n429_ = new_n426_ & ~new_n427_;
  assign \f[6]  = ~new_n428_ & ~new_n429_;
  assign new_n431_ = ~\a[7]  & ~\b[7] ;
  assign new_n432_ = \a[7]  & \b[7] ;
  assign new_n433_ = ~new_n431_ & ~new_n432_;
  assign new_n434_ = ~new_n425_ & ~new_n429_;
  assign new_n435_ = ~new_n433_ & new_n434_;
  assign new_n436_ = new_n433_ & ~new_n434_;
  assign \f[7]  = ~new_n435_ & ~new_n436_;
  assign new_n438_ = ~\a[8]  & ~\b[8] ;
  assign new_n439_ = \a[8]  & \b[8] ;
  assign new_n440_ = ~new_n438_ & ~new_n439_;
  assign new_n441_ = ~new_n432_ & ~new_n436_;
  assign new_n442_ = ~new_n440_ & new_n441_;
  assign new_n443_ = new_n440_ & ~new_n441_;
  assign \f[8]  = ~new_n442_ & ~new_n443_;
  assign new_n445_ = ~\a[9]  & ~\b[9] ;
  assign new_n446_ = \a[9]  & \b[9] ;
  assign new_n447_ = ~new_n445_ & ~new_n446_;
  assign new_n448_ = ~new_n439_ & ~new_n443_;
  assign new_n449_ = ~new_n447_ & new_n448_;
  assign new_n450_ = new_n447_ & ~new_n448_;
  assign \f[9]  = ~new_n449_ & ~new_n450_;
  assign new_n452_ = ~\a[10]  & ~\b[10] ;
  assign new_n453_ = \a[10]  & \b[10] ;
  assign new_n454_ = ~new_n452_ & ~new_n453_;
  assign new_n455_ = ~new_n446_ & ~new_n450_;
  assign new_n456_ = ~new_n454_ & new_n455_;
  assign new_n457_ = new_n454_ & ~new_n455_;
  assign \f[10]  = ~new_n456_ & ~new_n457_;
  assign new_n459_ = ~\a[11]  & ~\b[11] ;
  assign new_n460_ = \a[11]  & \b[11] ;
  assign new_n461_ = ~new_n459_ & ~new_n460_;
  assign new_n462_ = ~new_n453_ & ~new_n457_;
  assign new_n463_ = ~new_n461_ & new_n462_;
  assign new_n464_ = new_n461_ & ~new_n462_;
  assign \f[11]  = ~new_n463_ & ~new_n464_;
  assign new_n466_ = ~\a[12]  & ~\b[12] ;
  assign new_n467_ = \a[12]  & \b[12] ;
  assign new_n468_ = ~new_n466_ & ~new_n467_;
  assign new_n469_ = ~new_n460_ & ~new_n464_;
  assign new_n470_ = ~new_n468_ & new_n469_;
  assign new_n471_ = new_n468_ & ~new_n469_;
  assign \f[12]  = ~new_n470_ & ~new_n471_;
  assign new_n473_ = ~\a[13]  & ~\b[13] ;
  assign new_n474_ = \a[13]  & \b[13] ;
  assign new_n475_ = ~new_n473_ & ~new_n474_;
  assign new_n476_ = ~new_n467_ & ~new_n471_;
  assign new_n477_ = ~new_n475_ & new_n476_;
  assign new_n478_ = new_n475_ & ~new_n476_;
  assign \f[13]  = ~new_n477_ & ~new_n478_;
  assign new_n480_ = ~\a[14]  & ~\b[14] ;
  assign new_n481_ = \a[14]  & \b[14] ;
  assign new_n482_ = ~new_n480_ & ~new_n481_;
  assign new_n483_ = ~new_n474_ & ~new_n478_;
  assign new_n484_ = ~new_n482_ & new_n483_;
  assign new_n485_ = new_n482_ & ~new_n483_;
  assign \f[14]  = ~new_n484_ & ~new_n485_;
  assign new_n487_ = ~\a[15]  & ~\b[15] ;
  assign new_n488_ = \a[15]  & \b[15] ;
  assign new_n489_ = ~new_n487_ & ~new_n488_;
  assign new_n490_ = ~new_n481_ & ~new_n485_;
  assign new_n491_ = ~new_n489_ & new_n490_;
  assign new_n492_ = new_n489_ & ~new_n490_;
  assign \f[15]  = ~new_n491_ & ~new_n492_;
  assign new_n494_ = ~\a[16]  & ~\b[16] ;
  assign new_n495_ = \a[16]  & \b[16] ;
  assign new_n496_ = ~new_n494_ & ~new_n495_;
  assign new_n497_ = ~new_n488_ & ~new_n492_;
  assign new_n498_ = ~new_n496_ & new_n497_;
  assign new_n499_ = new_n496_ & ~new_n497_;
  assign \f[16]  = ~new_n498_ & ~new_n499_;
  assign new_n501_ = ~\a[17]  & ~\b[17] ;
  assign new_n502_ = \a[17]  & \b[17] ;
  assign new_n503_ = ~new_n501_ & ~new_n502_;
  assign new_n504_ = ~new_n495_ & ~new_n499_;
  assign new_n505_ = ~new_n503_ & new_n504_;
  assign new_n506_ = new_n503_ & ~new_n504_;
  assign \f[17]  = ~new_n505_ & ~new_n506_;
  assign new_n508_ = ~\a[18]  & ~\b[18] ;
  assign new_n509_ = \a[18]  & \b[18] ;
  assign new_n510_ = ~new_n508_ & ~new_n509_;
  assign new_n511_ = ~new_n502_ & ~new_n506_;
  assign new_n512_ = ~new_n510_ & new_n511_;
  assign new_n513_ = new_n510_ & ~new_n511_;
  assign \f[18]  = ~new_n512_ & ~new_n513_;
  assign new_n515_ = ~\a[19]  & ~\b[19] ;
  assign new_n516_ = \a[19]  & \b[19] ;
  assign new_n517_ = ~new_n515_ & ~new_n516_;
  assign new_n518_ = ~new_n509_ & ~new_n513_;
  assign new_n519_ = ~new_n517_ & new_n518_;
  assign new_n520_ = new_n517_ & ~new_n518_;
  assign \f[19]  = ~new_n519_ & ~new_n520_;
  assign new_n522_ = ~\a[20]  & ~\b[20] ;
  assign new_n523_ = \a[20]  & \b[20] ;
  assign new_n524_ = ~new_n522_ & ~new_n523_;
  assign new_n525_ = ~new_n516_ & ~new_n520_;
  assign new_n526_ = ~new_n524_ & new_n525_;
  assign new_n527_ = new_n524_ & ~new_n525_;
  assign \f[20]  = ~new_n526_ & ~new_n527_;
  assign new_n529_ = ~\a[21]  & ~\b[21] ;
  assign new_n530_ = \a[21]  & \b[21] ;
  assign new_n531_ = ~new_n529_ & ~new_n530_;
  assign new_n532_ = ~new_n523_ & ~new_n527_;
  assign new_n533_ = ~new_n531_ & new_n532_;
  assign new_n534_ = new_n531_ & ~new_n532_;
  assign \f[21]  = ~new_n533_ & ~new_n534_;
  assign new_n536_ = ~\a[22]  & ~\b[22] ;
  assign new_n537_ = \a[22]  & \b[22] ;
  assign new_n538_ = ~new_n536_ & ~new_n537_;
  assign new_n539_ = ~new_n530_ & ~new_n534_;
  assign new_n540_ = ~new_n538_ & new_n539_;
  assign new_n541_ = new_n538_ & ~new_n539_;
  assign \f[22]  = ~new_n540_ & ~new_n541_;
  assign new_n543_ = ~\a[23]  & ~\b[23] ;
  assign new_n544_ = \a[23]  & \b[23] ;
  assign new_n545_ = ~new_n543_ & ~new_n544_;
  assign new_n546_ = ~new_n537_ & ~new_n541_;
  assign new_n547_ = ~new_n545_ & new_n546_;
  assign new_n548_ = new_n545_ & ~new_n546_;
  assign \f[23]  = ~new_n547_ & ~new_n548_;
  assign new_n550_ = ~\a[24]  & ~\b[24] ;
  assign new_n551_ = \a[24]  & \b[24] ;
  assign new_n552_ = ~new_n550_ & ~new_n551_;
  assign new_n553_ = ~new_n544_ & ~new_n548_;
  assign new_n554_ = ~new_n552_ & new_n553_;
  assign new_n555_ = new_n552_ & ~new_n553_;
  assign \f[24]  = ~new_n554_ & ~new_n555_;
  assign new_n557_ = ~\a[25]  & ~\b[25] ;
  assign new_n558_ = \a[25]  & \b[25] ;
  assign new_n559_ = ~new_n557_ & ~new_n558_;
  assign new_n560_ = ~new_n551_ & ~new_n555_;
  assign new_n561_ = ~new_n559_ & new_n560_;
  assign new_n562_ = new_n559_ & ~new_n560_;
  assign \f[25]  = ~new_n561_ & ~new_n562_;
  assign new_n564_ = ~\a[26]  & ~\b[26] ;
  assign new_n565_ = \a[26]  & \b[26] ;
  assign new_n566_ = ~new_n564_ & ~new_n565_;
  assign new_n567_ = ~new_n558_ & ~new_n562_;
  assign new_n568_ = ~new_n566_ & new_n567_;
  assign new_n569_ = new_n566_ & ~new_n567_;
  assign \f[26]  = ~new_n568_ & ~new_n569_;
  assign new_n571_ = ~\a[27]  & ~\b[27] ;
  assign new_n572_ = \a[27]  & \b[27] ;
  assign new_n573_ = ~new_n571_ & ~new_n572_;
  assign new_n574_ = ~new_n565_ & ~new_n569_;
  assign new_n575_ = ~new_n573_ & new_n574_;
  assign new_n576_ = new_n573_ & ~new_n574_;
  assign \f[27]  = ~new_n575_ & ~new_n576_;
  assign new_n578_ = ~\a[28]  & ~\b[28] ;
  assign new_n579_ = \a[28]  & \b[28] ;
  assign new_n580_ = ~new_n578_ & ~new_n579_;
  assign new_n581_ = ~new_n572_ & ~new_n576_;
  assign new_n582_ = ~new_n580_ & new_n581_;
  assign new_n583_ = new_n580_ & ~new_n581_;
  assign \f[28]  = ~new_n582_ & ~new_n583_;
  assign new_n585_ = ~\a[29]  & ~\b[29] ;
  assign new_n586_ = \a[29]  & \b[29] ;
  assign new_n587_ = ~new_n585_ & ~new_n586_;
  assign new_n588_ = ~new_n579_ & ~new_n583_;
  assign new_n589_ = ~new_n587_ & new_n588_;
  assign new_n590_ = new_n587_ & ~new_n588_;
  assign \f[29]  = ~new_n589_ & ~new_n590_;
  assign new_n592_ = ~\a[30]  & ~\b[30] ;
  assign new_n593_ = \a[30]  & \b[30] ;
  assign new_n594_ = ~new_n592_ & ~new_n593_;
  assign new_n595_ = ~new_n586_ & ~new_n590_;
  assign new_n596_ = ~new_n594_ & new_n595_;
  assign new_n597_ = new_n594_ & ~new_n595_;
  assign \f[30]  = ~new_n596_ & ~new_n597_;
  assign new_n599_ = ~\a[31]  & ~\b[31] ;
  assign new_n600_ = \a[31]  & \b[31] ;
  assign new_n601_ = ~new_n599_ & ~new_n600_;
  assign new_n602_ = ~new_n593_ & ~new_n597_;
  assign new_n603_ = ~new_n601_ & new_n602_;
  assign new_n604_ = new_n601_ & ~new_n602_;
  assign \f[31]  = ~new_n603_ & ~new_n604_;
  assign new_n606_ = ~\a[32]  & ~\b[32] ;
  assign new_n607_ = \a[32]  & \b[32] ;
  assign new_n608_ = ~new_n606_ & ~new_n607_;
  assign new_n609_ = ~new_n600_ & ~new_n604_;
  assign new_n610_ = ~new_n608_ & new_n609_;
  assign new_n611_ = new_n608_ & ~new_n609_;
  assign \f[32]  = ~new_n610_ & ~new_n611_;
  assign new_n613_ = ~\a[33]  & ~\b[33] ;
  assign new_n614_ = \a[33]  & \b[33] ;
  assign new_n615_ = ~new_n613_ & ~new_n614_;
  assign new_n616_ = ~new_n607_ & ~new_n611_;
  assign new_n617_ = ~new_n615_ & new_n616_;
  assign new_n618_ = new_n615_ & ~new_n616_;
  assign \f[33]  = ~new_n617_ & ~new_n618_;
  assign new_n620_ = ~\a[34]  & ~\b[34] ;
  assign new_n621_ = \a[34]  & \b[34] ;
  assign new_n622_ = ~new_n620_ & ~new_n621_;
  assign new_n623_ = ~new_n614_ & ~new_n618_;
  assign new_n624_ = ~new_n622_ & new_n623_;
  assign new_n625_ = new_n622_ & ~new_n623_;
  assign \f[34]  = ~new_n624_ & ~new_n625_;
  assign new_n627_ = ~\a[35]  & ~\b[35] ;
  assign new_n628_ = \a[35]  & \b[35] ;
  assign new_n629_ = ~new_n627_ & ~new_n628_;
  assign new_n630_ = ~new_n621_ & ~new_n625_;
  assign new_n631_ = ~new_n629_ & new_n630_;
  assign new_n632_ = new_n629_ & ~new_n630_;
  assign \f[35]  = ~new_n631_ & ~new_n632_;
  assign new_n634_ = ~\a[36]  & ~\b[36] ;
  assign new_n635_ = \a[36]  & \b[36] ;
  assign new_n636_ = ~new_n634_ & ~new_n635_;
  assign new_n637_ = ~new_n628_ & ~new_n632_;
  assign new_n638_ = ~new_n636_ & new_n637_;
  assign new_n639_ = new_n636_ & ~new_n637_;
  assign \f[36]  = ~new_n638_ & ~new_n639_;
  assign new_n641_ = ~\a[37]  & ~\b[37] ;
  assign new_n642_ = \a[37]  & \b[37] ;
  assign new_n643_ = ~new_n641_ & ~new_n642_;
  assign new_n644_ = ~new_n635_ & ~new_n639_;
  assign new_n645_ = ~new_n643_ & new_n644_;
  assign new_n646_ = new_n643_ & ~new_n644_;
  assign \f[37]  = ~new_n645_ & ~new_n646_;
  assign new_n648_ = ~\a[38]  & ~\b[38] ;
  assign new_n649_ = \a[38]  & \b[38] ;
  assign new_n650_ = ~new_n648_ & ~new_n649_;
  assign new_n651_ = ~new_n642_ & ~new_n646_;
  assign new_n652_ = ~new_n650_ & new_n651_;
  assign new_n653_ = new_n650_ & ~new_n651_;
  assign \f[38]  = ~new_n652_ & ~new_n653_;
  assign new_n655_ = ~\a[39]  & ~\b[39] ;
  assign new_n656_ = \a[39]  & \b[39] ;
  assign new_n657_ = ~new_n655_ & ~new_n656_;
  assign new_n658_ = ~new_n649_ & ~new_n653_;
  assign new_n659_ = ~new_n657_ & new_n658_;
  assign new_n660_ = new_n657_ & ~new_n658_;
  assign \f[39]  = ~new_n659_ & ~new_n660_;
  assign new_n662_ = ~\a[40]  & ~\b[40] ;
  assign new_n663_ = \a[40]  & \b[40] ;
  assign new_n664_ = ~new_n662_ & ~new_n663_;
  assign new_n665_ = ~new_n656_ & ~new_n660_;
  assign new_n666_ = ~new_n664_ & new_n665_;
  assign new_n667_ = new_n664_ & ~new_n665_;
  assign \f[40]  = ~new_n666_ & ~new_n667_;
  assign new_n669_ = ~\a[41]  & ~\b[41] ;
  assign new_n670_ = \a[41]  & \b[41] ;
  assign new_n671_ = ~new_n669_ & ~new_n670_;
  assign new_n672_ = ~new_n663_ & ~new_n667_;
  assign new_n673_ = ~new_n671_ & new_n672_;
  assign new_n674_ = new_n671_ & ~new_n672_;
  assign \f[41]  = ~new_n673_ & ~new_n674_;
  assign new_n676_ = ~\a[42]  & ~\b[42] ;
  assign new_n677_ = \a[42]  & \b[42] ;
  assign new_n678_ = ~new_n676_ & ~new_n677_;
  assign new_n679_ = ~new_n670_ & ~new_n674_;
  assign new_n680_ = ~new_n678_ & new_n679_;
  assign new_n681_ = new_n678_ & ~new_n679_;
  assign \f[42]  = ~new_n680_ & ~new_n681_;
  assign new_n683_ = ~\a[43]  & ~\b[43] ;
  assign new_n684_ = \a[43]  & \b[43] ;
  assign new_n685_ = ~new_n683_ & ~new_n684_;
  assign new_n686_ = ~new_n677_ & ~new_n681_;
  assign new_n687_ = ~new_n685_ & new_n686_;
  assign new_n688_ = new_n685_ & ~new_n686_;
  assign \f[43]  = ~new_n687_ & ~new_n688_;
  assign new_n690_ = ~\a[44]  & ~\b[44] ;
  assign new_n691_ = \a[44]  & \b[44] ;
  assign new_n692_ = ~new_n690_ & ~new_n691_;
  assign new_n693_ = ~new_n684_ & ~new_n688_;
  assign new_n694_ = ~new_n692_ & new_n693_;
  assign new_n695_ = new_n692_ & ~new_n693_;
  assign \f[44]  = ~new_n694_ & ~new_n695_;
  assign new_n697_ = ~\a[45]  & ~\b[45] ;
  assign new_n698_ = \a[45]  & \b[45] ;
  assign new_n699_ = ~new_n697_ & ~new_n698_;
  assign new_n700_ = ~new_n691_ & ~new_n695_;
  assign new_n701_ = ~new_n699_ & new_n700_;
  assign new_n702_ = new_n699_ & ~new_n700_;
  assign \f[45]  = ~new_n701_ & ~new_n702_;
  assign new_n704_ = ~\a[46]  & ~\b[46] ;
  assign new_n705_ = \a[46]  & \b[46] ;
  assign new_n706_ = ~new_n704_ & ~new_n705_;
  assign new_n707_ = ~new_n698_ & ~new_n702_;
  assign new_n708_ = ~new_n706_ & new_n707_;
  assign new_n709_ = new_n706_ & ~new_n707_;
  assign \f[46]  = ~new_n708_ & ~new_n709_;
  assign new_n711_ = ~\a[47]  & ~\b[47] ;
  assign new_n712_ = \a[47]  & \b[47] ;
  assign new_n713_ = ~new_n711_ & ~new_n712_;
  assign new_n714_ = ~new_n705_ & ~new_n709_;
  assign new_n715_ = ~new_n713_ & new_n714_;
  assign new_n716_ = new_n713_ & ~new_n714_;
  assign \f[47]  = ~new_n715_ & ~new_n716_;
  assign new_n718_ = ~\a[48]  & ~\b[48] ;
  assign new_n719_ = \a[48]  & \b[48] ;
  assign new_n720_ = ~new_n718_ & ~new_n719_;
  assign new_n721_ = ~new_n712_ & ~new_n716_;
  assign new_n722_ = ~new_n720_ & new_n721_;
  assign new_n723_ = new_n720_ & ~new_n721_;
  assign \f[48]  = ~new_n722_ & ~new_n723_;
  assign new_n725_ = ~\a[49]  & ~\b[49] ;
  assign new_n726_ = \a[49]  & \b[49] ;
  assign new_n727_ = ~new_n725_ & ~new_n726_;
  assign new_n728_ = ~new_n719_ & ~new_n723_;
  assign new_n729_ = ~new_n727_ & new_n728_;
  assign new_n730_ = new_n727_ & ~new_n728_;
  assign \f[49]  = ~new_n729_ & ~new_n730_;
  assign new_n732_ = ~\a[50]  & ~\b[50] ;
  assign new_n733_ = \a[50]  & \b[50] ;
  assign new_n734_ = ~new_n732_ & ~new_n733_;
  assign new_n735_ = ~new_n726_ & ~new_n730_;
  assign new_n736_ = ~new_n734_ & new_n735_;
  assign new_n737_ = new_n734_ & ~new_n735_;
  assign \f[50]  = ~new_n736_ & ~new_n737_;
  assign new_n739_ = ~\a[51]  & ~\b[51] ;
  assign new_n740_ = \a[51]  & \b[51] ;
  assign new_n741_ = ~new_n739_ & ~new_n740_;
  assign new_n742_ = ~new_n733_ & ~new_n737_;
  assign new_n743_ = ~new_n741_ & new_n742_;
  assign new_n744_ = new_n741_ & ~new_n742_;
  assign \f[51]  = ~new_n743_ & ~new_n744_;
  assign new_n746_ = ~\a[52]  & ~\b[52] ;
  assign new_n747_ = \a[52]  & \b[52] ;
  assign new_n748_ = ~new_n746_ & ~new_n747_;
  assign new_n749_ = ~new_n740_ & ~new_n744_;
  assign new_n750_ = ~new_n748_ & new_n749_;
  assign new_n751_ = new_n748_ & ~new_n749_;
  assign \f[52]  = ~new_n750_ & ~new_n751_;
  assign new_n753_ = ~\a[53]  & ~\b[53] ;
  assign new_n754_ = \a[53]  & \b[53] ;
  assign new_n755_ = ~new_n753_ & ~new_n754_;
  assign new_n756_ = ~new_n747_ & ~new_n751_;
  assign new_n757_ = ~new_n755_ & new_n756_;
  assign new_n758_ = new_n755_ & ~new_n756_;
  assign \f[53]  = ~new_n757_ & ~new_n758_;
  assign new_n760_ = ~\a[54]  & ~\b[54] ;
  assign new_n761_ = \a[54]  & \b[54] ;
  assign new_n762_ = ~new_n760_ & ~new_n761_;
  assign new_n763_ = ~new_n754_ & ~new_n758_;
  assign new_n764_ = ~new_n762_ & new_n763_;
  assign new_n765_ = new_n762_ & ~new_n763_;
  assign \f[54]  = ~new_n764_ & ~new_n765_;
  assign new_n767_ = ~\a[55]  & ~\b[55] ;
  assign new_n768_ = \a[55]  & \b[55] ;
  assign new_n769_ = ~new_n767_ & ~new_n768_;
  assign new_n770_ = ~new_n761_ & ~new_n765_;
  assign new_n771_ = ~new_n769_ & new_n770_;
  assign new_n772_ = new_n769_ & ~new_n770_;
  assign \f[55]  = ~new_n771_ & ~new_n772_;
  assign new_n774_ = ~\a[56]  & ~\b[56] ;
  assign new_n775_ = \a[56]  & \b[56] ;
  assign new_n776_ = ~new_n774_ & ~new_n775_;
  assign new_n777_ = ~new_n768_ & ~new_n772_;
  assign new_n778_ = ~new_n776_ & new_n777_;
  assign new_n779_ = new_n776_ & ~new_n777_;
  assign \f[56]  = ~new_n778_ & ~new_n779_;
  assign new_n781_ = ~\a[57]  & ~\b[57] ;
  assign new_n782_ = \a[57]  & \b[57] ;
  assign new_n783_ = ~new_n781_ & ~new_n782_;
  assign new_n784_ = ~new_n775_ & ~new_n779_;
  assign new_n785_ = ~new_n783_ & new_n784_;
  assign new_n786_ = new_n783_ & ~new_n784_;
  assign \f[57]  = ~new_n785_ & ~new_n786_;
  assign new_n788_ = ~\a[58]  & ~\b[58] ;
  assign new_n789_ = \a[58]  & \b[58] ;
  assign new_n790_ = ~new_n788_ & ~new_n789_;
  assign new_n791_ = ~new_n782_ & ~new_n786_;
  assign new_n792_ = ~new_n790_ & new_n791_;
  assign new_n793_ = new_n790_ & ~new_n791_;
  assign \f[58]  = ~new_n792_ & ~new_n793_;
  assign new_n795_ = ~\a[59]  & ~\b[59] ;
  assign new_n796_ = \a[59]  & \b[59] ;
  assign new_n797_ = ~new_n795_ & ~new_n796_;
  assign new_n798_ = ~new_n789_ & ~new_n793_;
  assign new_n799_ = ~new_n797_ & new_n798_;
  assign new_n800_ = new_n797_ & ~new_n798_;
  assign \f[59]  = ~new_n799_ & ~new_n800_;
  assign new_n802_ = ~\a[60]  & ~\b[60] ;
  assign new_n803_ = \a[60]  & \b[60] ;
  assign new_n804_ = ~new_n802_ & ~new_n803_;
  assign new_n805_ = ~new_n796_ & ~new_n800_;
  assign new_n806_ = ~new_n804_ & new_n805_;
  assign new_n807_ = new_n804_ & ~new_n805_;
  assign \f[60]  = ~new_n806_ & ~new_n807_;
  assign new_n809_ = ~\a[61]  & ~\b[61] ;
  assign new_n810_ = \a[61]  & \b[61] ;
  assign new_n811_ = ~new_n809_ & ~new_n810_;
  assign new_n812_ = ~new_n803_ & ~new_n807_;
  assign new_n813_ = ~new_n811_ & new_n812_;
  assign new_n814_ = new_n811_ & ~new_n812_;
  assign \f[61]  = ~new_n813_ & ~new_n814_;
  assign new_n816_ = ~\a[62]  & ~\b[62] ;
  assign new_n817_ = \a[62]  & \b[62] ;
  assign new_n818_ = ~new_n816_ & ~new_n817_;
  assign new_n819_ = ~new_n810_ & ~new_n814_;
  assign new_n820_ = ~new_n818_ & new_n819_;
  assign new_n821_ = new_n818_ & ~new_n819_;
  assign \f[62]  = ~new_n820_ & ~new_n821_;
  assign new_n823_ = ~\a[63]  & ~\b[63] ;
  assign new_n824_ = \a[63]  & \b[63] ;
  assign new_n825_ = ~new_n823_ & ~new_n824_;
  assign new_n826_ = ~new_n817_ & ~new_n821_;
  assign new_n827_ = ~new_n825_ & new_n826_;
  assign new_n828_ = new_n825_ & ~new_n826_;
  assign \f[63]  = ~new_n827_ & ~new_n828_;
  assign new_n830_ = ~\a[64]  & ~\b[64] ;
  assign new_n831_ = \a[64]  & \b[64] ;
  assign new_n832_ = ~new_n830_ & ~new_n831_;
  assign new_n833_ = ~new_n824_ & ~new_n828_;
  assign new_n834_ = ~new_n832_ & new_n833_;
  assign new_n835_ = new_n832_ & ~new_n833_;
  assign \f[64]  = ~new_n834_ & ~new_n835_;
  assign new_n837_ = ~\a[65]  & ~\b[65] ;
  assign new_n838_ = \a[65]  & \b[65] ;
  assign new_n839_ = ~new_n837_ & ~new_n838_;
  assign new_n840_ = ~new_n831_ & ~new_n835_;
  assign new_n841_ = ~new_n839_ & new_n840_;
  assign new_n842_ = new_n839_ & ~new_n840_;
  assign \f[65]  = ~new_n841_ & ~new_n842_;
  assign new_n844_ = ~\a[66]  & ~\b[66] ;
  assign new_n845_ = \a[66]  & \b[66] ;
  assign new_n846_ = ~new_n844_ & ~new_n845_;
  assign new_n847_ = ~new_n838_ & ~new_n842_;
  assign new_n848_ = ~new_n846_ & new_n847_;
  assign new_n849_ = new_n846_ & ~new_n847_;
  assign \f[66]  = ~new_n848_ & ~new_n849_;
  assign new_n851_ = ~\a[67]  & ~\b[67] ;
  assign new_n852_ = \a[67]  & \b[67] ;
  assign new_n853_ = ~new_n851_ & ~new_n852_;
  assign new_n854_ = ~new_n845_ & ~new_n849_;
  assign new_n855_ = ~new_n853_ & new_n854_;
  assign new_n856_ = new_n853_ & ~new_n854_;
  assign \f[67]  = ~new_n855_ & ~new_n856_;
  assign new_n858_ = ~\a[68]  & ~\b[68] ;
  assign new_n859_ = \a[68]  & \b[68] ;
  assign new_n860_ = ~new_n858_ & ~new_n859_;
  assign new_n861_ = ~new_n852_ & ~new_n856_;
  assign new_n862_ = ~new_n860_ & new_n861_;
  assign new_n863_ = new_n860_ & ~new_n861_;
  assign \f[68]  = ~new_n862_ & ~new_n863_;
  assign new_n865_ = ~\a[69]  & ~\b[69] ;
  assign new_n866_ = \a[69]  & \b[69] ;
  assign new_n867_ = ~new_n865_ & ~new_n866_;
  assign new_n868_ = ~new_n859_ & ~new_n863_;
  assign new_n869_ = ~new_n867_ & new_n868_;
  assign new_n870_ = new_n867_ & ~new_n868_;
  assign \f[69]  = ~new_n869_ & ~new_n870_;
  assign new_n872_ = ~\a[70]  & ~\b[70] ;
  assign new_n873_ = \a[70]  & \b[70] ;
  assign new_n874_ = ~new_n872_ & ~new_n873_;
  assign new_n875_ = ~new_n866_ & ~new_n870_;
  assign new_n876_ = ~new_n874_ & new_n875_;
  assign new_n877_ = new_n874_ & ~new_n875_;
  assign \f[70]  = ~new_n876_ & ~new_n877_;
  assign new_n879_ = ~\a[71]  & ~\b[71] ;
  assign new_n880_ = \a[71]  & \b[71] ;
  assign new_n881_ = ~new_n879_ & ~new_n880_;
  assign new_n882_ = ~new_n873_ & ~new_n877_;
  assign new_n883_ = ~new_n881_ & new_n882_;
  assign new_n884_ = new_n881_ & ~new_n882_;
  assign \f[71]  = ~new_n883_ & ~new_n884_;
  assign new_n886_ = ~\a[72]  & ~\b[72] ;
  assign new_n887_ = \a[72]  & \b[72] ;
  assign new_n888_ = ~new_n886_ & ~new_n887_;
  assign new_n889_ = ~new_n880_ & ~new_n884_;
  assign new_n890_ = ~new_n888_ & new_n889_;
  assign new_n891_ = new_n888_ & ~new_n889_;
  assign \f[72]  = ~new_n890_ & ~new_n891_;
  assign new_n893_ = ~\a[73]  & ~\b[73] ;
  assign new_n894_ = \a[73]  & \b[73] ;
  assign new_n895_ = ~new_n893_ & ~new_n894_;
  assign new_n896_ = ~new_n887_ & ~new_n891_;
  assign new_n897_ = ~new_n895_ & new_n896_;
  assign new_n898_ = new_n895_ & ~new_n896_;
  assign \f[73]  = ~new_n897_ & ~new_n898_;
  assign new_n900_ = ~\a[74]  & ~\b[74] ;
  assign new_n901_ = \a[74]  & \b[74] ;
  assign new_n902_ = ~new_n900_ & ~new_n901_;
  assign new_n903_ = ~new_n894_ & ~new_n898_;
  assign new_n904_ = ~new_n902_ & new_n903_;
  assign new_n905_ = new_n902_ & ~new_n903_;
  assign \f[74]  = ~new_n904_ & ~new_n905_;
  assign new_n907_ = ~\a[75]  & ~\b[75] ;
  assign new_n908_ = \a[75]  & \b[75] ;
  assign new_n909_ = ~new_n907_ & ~new_n908_;
  assign new_n910_ = ~new_n901_ & ~new_n905_;
  assign new_n911_ = ~new_n909_ & new_n910_;
  assign new_n912_ = new_n909_ & ~new_n910_;
  assign \f[75]  = ~new_n911_ & ~new_n912_;
  assign new_n914_ = ~\a[76]  & ~\b[76] ;
  assign new_n915_ = \a[76]  & \b[76] ;
  assign new_n916_ = ~new_n914_ & ~new_n915_;
  assign new_n917_ = ~new_n908_ & ~new_n912_;
  assign new_n918_ = ~new_n916_ & new_n917_;
  assign new_n919_ = new_n916_ & ~new_n917_;
  assign \f[76]  = ~new_n918_ & ~new_n919_;
  assign new_n921_ = ~\a[77]  & ~\b[77] ;
  assign new_n922_ = \a[77]  & \b[77] ;
  assign new_n923_ = ~new_n921_ & ~new_n922_;
  assign new_n924_ = ~new_n915_ & ~new_n919_;
  assign new_n925_ = ~new_n923_ & new_n924_;
  assign new_n926_ = new_n923_ & ~new_n924_;
  assign \f[77]  = ~new_n925_ & ~new_n926_;
  assign new_n928_ = ~\a[78]  & ~\b[78] ;
  assign new_n929_ = \a[78]  & \b[78] ;
  assign new_n930_ = ~new_n928_ & ~new_n929_;
  assign new_n931_ = ~new_n922_ & ~new_n926_;
  assign new_n932_ = ~new_n930_ & new_n931_;
  assign new_n933_ = new_n930_ & ~new_n931_;
  assign \f[78]  = ~new_n932_ & ~new_n933_;
  assign new_n935_ = ~\a[79]  & ~\b[79] ;
  assign new_n936_ = \a[79]  & \b[79] ;
  assign new_n937_ = ~new_n935_ & ~new_n936_;
  assign new_n938_ = ~new_n929_ & ~new_n933_;
  assign new_n939_ = ~new_n937_ & new_n938_;
  assign new_n940_ = new_n937_ & ~new_n938_;
  assign \f[79]  = ~new_n939_ & ~new_n940_;
  assign new_n942_ = ~\a[80]  & ~\b[80] ;
  assign new_n943_ = \a[80]  & \b[80] ;
  assign new_n944_ = ~new_n942_ & ~new_n943_;
  assign new_n945_ = ~new_n936_ & ~new_n940_;
  assign new_n946_ = ~new_n944_ & new_n945_;
  assign new_n947_ = new_n944_ & ~new_n945_;
  assign \f[80]  = ~new_n946_ & ~new_n947_;
  assign new_n949_ = ~\a[81]  & ~\b[81] ;
  assign new_n950_ = \a[81]  & \b[81] ;
  assign new_n951_ = ~new_n949_ & ~new_n950_;
  assign new_n952_ = ~new_n943_ & ~new_n947_;
  assign new_n953_ = ~new_n951_ & new_n952_;
  assign new_n954_ = new_n951_ & ~new_n952_;
  assign \f[81]  = ~new_n953_ & ~new_n954_;
  assign new_n956_ = ~\a[82]  & ~\b[82] ;
  assign new_n957_ = \a[82]  & \b[82] ;
  assign new_n958_ = ~new_n956_ & ~new_n957_;
  assign new_n959_ = ~new_n950_ & ~new_n954_;
  assign new_n960_ = ~new_n958_ & new_n959_;
  assign new_n961_ = new_n958_ & ~new_n959_;
  assign \f[82]  = ~new_n960_ & ~new_n961_;
  assign new_n963_ = ~\a[83]  & ~\b[83] ;
  assign new_n964_ = \a[83]  & \b[83] ;
  assign new_n965_ = ~new_n963_ & ~new_n964_;
  assign new_n966_ = ~new_n957_ & ~new_n961_;
  assign new_n967_ = ~new_n965_ & new_n966_;
  assign new_n968_ = new_n965_ & ~new_n966_;
  assign \f[83]  = ~new_n967_ & ~new_n968_;
  assign new_n970_ = ~\a[84]  & ~\b[84] ;
  assign new_n971_ = \a[84]  & \b[84] ;
  assign new_n972_ = ~new_n970_ & ~new_n971_;
  assign new_n973_ = ~new_n964_ & ~new_n968_;
  assign new_n974_ = ~new_n972_ & new_n973_;
  assign new_n975_ = new_n972_ & ~new_n973_;
  assign \f[84]  = ~new_n974_ & ~new_n975_;
  assign new_n977_ = ~\a[85]  & ~\b[85] ;
  assign new_n978_ = \a[85]  & \b[85] ;
  assign new_n979_ = ~new_n977_ & ~new_n978_;
  assign new_n980_ = ~new_n971_ & ~new_n975_;
  assign new_n981_ = ~new_n979_ & new_n980_;
  assign new_n982_ = new_n979_ & ~new_n980_;
  assign \f[85]  = ~new_n981_ & ~new_n982_;
  assign new_n984_ = ~\a[86]  & ~\b[86] ;
  assign new_n985_ = \a[86]  & \b[86] ;
  assign new_n986_ = ~new_n984_ & ~new_n985_;
  assign new_n987_ = ~new_n978_ & ~new_n982_;
  assign new_n988_ = ~new_n986_ & new_n987_;
  assign new_n989_ = new_n986_ & ~new_n987_;
  assign \f[86]  = ~new_n988_ & ~new_n989_;
  assign new_n991_ = ~\a[87]  & ~\b[87] ;
  assign new_n992_ = \a[87]  & \b[87] ;
  assign new_n993_ = ~new_n991_ & ~new_n992_;
  assign new_n994_ = ~new_n985_ & ~new_n989_;
  assign new_n995_ = ~new_n993_ & new_n994_;
  assign new_n996_ = new_n993_ & ~new_n994_;
  assign \f[87]  = ~new_n995_ & ~new_n996_;
  assign new_n998_ = ~\a[88]  & ~\b[88] ;
  assign new_n999_ = \a[88]  & \b[88] ;
  assign new_n1000_ = ~new_n998_ & ~new_n999_;
  assign new_n1001_ = ~new_n992_ & ~new_n996_;
  assign new_n1002_ = ~new_n1000_ & new_n1001_;
  assign new_n1003_ = new_n1000_ & ~new_n1001_;
  assign \f[88]  = ~new_n1002_ & ~new_n1003_;
  assign new_n1005_ = ~\a[89]  & ~\b[89] ;
  assign new_n1006_ = \a[89]  & \b[89] ;
  assign new_n1007_ = ~new_n1005_ & ~new_n1006_;
  assign new_n1008_ = ~new_n999_ & ~new_n1003_;
  assign new_n1009_ = ~new_n1007_ & new_n1008_;
  assign new_n1010_ = new_n1007_ & ~new_n1008_;
  assign \f[89]  = ~new_n1009_ & ~new_n1010_;
  assign new_n1012_ = ~\a[90]  & ~\b[90] ;
  assign new_n1013_ = \a[90]  & \b[90] ;
  assign new_n1014_ = ~new_n1012_ & ~new_n1013_;
  assign new_n1015_ = ~new_n1006_ & ~new_n1010_;
  assign new_n1016_ = ~new_n1014_ & new_n1015_;
  assign new_n1017_ = new_n1014_ & ~new_n1015_;
  assign \f[90]  = ~new_n1016_ & ~new_n1017_;
  assign new_n1019_ = ~\a[91]  & ~\b[91] ;
  assign new_n1020_ = \a[91]  & \b[91] ;
  assign new_n1021_ = ~new_n1019_ & ~new_n1020_;
  assign new_n1022_ = ~new_n1013_ & ~new_n1017_;
  assign new_n1023_ = ~new_n1021_ & new_n1022_;
  assign new_n1024_ = new_n1021_ & ~new_n1022_;
  assign \f[91]  = ~new_n1023_ & ~new_n1024_;
  assign new_n1026_ = ~\a[92]  & ~\b[92] ;
  assign new_n1027_ = \a[92]  & \b[92] ;
  assign new_n1028_ = ~new_n1026_ & ~new_n1027_;
  assign new_n1029_ = ~new_n1020_ & ~new_n1024_;
  assign new_n1030_ = ~new_n1028_ & new_n1029_;
  assign new_n1031_ = new_n1028_ & ~new_n1029_;
  assign \f[92]  = ~new_n1030_ & ~new_n1031_;
  assign new_n1033_ = ~\a[93]  & ~\b[93] ;
  assign new_n1034_ = \a[93]  & \b[93] ;
  assign new_n1035_ = ~new_n1033_ & ~new_n1034_;
  assign new_n1036_ = ~new_n1027_ & ~new_n1031_;
  assign new_n1037_ = ~new_n1035_ & new_n1036_;
  assign new_n1038_ = new_n1035_ & ~new_n1036_;
  assign \f[93]  = ~new_n1037_ & ~new_n1038_;
  assign new_n1040_ = ~\a[94]  & ~\b[94] ;
  assign new_n1041_ = \a[94]  & \b[94] ;
  assign new_n1042_ = ~new_n1040_ & ~new_n1041_;
  assign new_n1043_ = ~new_n1034_ & ~new_n1038_;
  assign new_n1044_ = ~new_n1042_ & new_n1043_;
  assign new_n1045_ = new_n1042_ & ~new_n1043_;
  assign \f[94]  = ~new_n1044_ & ~new_n1045_;
  assign new_n1047_ = ~\a[95]  & ~\b[95] ;
  assign new_n1048_ = \a[95]  & \b[95] ;
  assign new_n1049_ = ~new_n1047_ & ~new_n1048_;
  assign new_n1050_ = ~new_n1041_ & ~new_n1045_;
  assign new_n1051_ = ~new_n1049_ & new_n1050_;
  assign new_n1052_ = new_n1049_ & ~new_n1050_;
  assign \f[95]  = ~new_n1051_ & ~new_n1052_;
  assign new_n1054_ = ~\a[96]  & ~\b[96] ;
  assign new_n1055_ = \a[96]  & \b[96] ;
  assign new_n1056_ = ~new_n1054_ & ~new_n1055_;
  assign new_n1057_ = ~new_n1048_ & ~new_n1052_;
  assign new_n1058_ = ~new_n1056_ & new_n1057_;
  assign new_n1059_ = new_n1056_ & ~new_n1057_;
  assign \f[96]  = ~new_n1058_ & ~new_n1059_;
  assign new_n1061_ = ~\a[97]  & ~\b[97] ;
  assign new_n1062_ = \a[97]  & \b[97] ;
  assign new_n1063_ = ~new_n1061_ & ~new_n1062_;
  assign new_n1064_ = ~new_n1055_ & ~new_n1059_;
  assign new_n1065_ = ~new_n1063_ & new_n1064_;
  assign new_n1066_ = new_n1063_ & ~new_n1064_;
  assign \f[97]  = ~new_n1065_ & ~new_n1066_;
  assign new_n1068_ = ~\a[98]  & ~\b[98] ;
  assign new_n1069_ = \a[98]  & \b[98] ;
  assign new_n1070_ = ~new_n1068_ & ~new_n1069_;
  assign new_n1071_ = ~new_n1062_ & ~new_n1066_;
  assign new_n1072_ = ~new_n1070_ & new_n1071_;
  assign new_n1073_ = new_n1070_ & ~new_n1071_;
  assign \f[98]  = ~new_n1072_ & ~new_n1073_;
  assign new_n1075_ = ~\a[99]  & ~\b[99] ;
  assign new_n1076_ = \a[99]  & \b[99] ;
  assign new_n1077_ = ~new_n1075_ & ~new_n1076_;
  assign new_n1078_ = ~new_n1069_ & ~new_n1073_;
  assign new_n1079_ = ~new_n1077_ & new_n1078_;
  assign new_n1080_ = new_n1077_ & ~new_n1078_;
  assign \f[99]  = ~new_n1079_ & ~new_n1080_;
  assign new_n1082_ = ~\a[100]  & ~\b[100] ;
  assign new_n1083_ = \a[100]  & \b[100] ;
  assign new_n1084_ = ~new_n1082_ & ~new_n1083_;
  assign new_n1085_ = ~new_n1076_ & ~new_n1080_;
  assign new_n1086_ = ~new_n1084_ & new_n1085_;
  assign new_n1087_ = new_n1084_ & ~new_n1085_;
  assign \f[100]  = ~new_n1086_ & ~new_n1087_;
  assign new_n1089_ = ~\a[101]  & ~\b[101] ;
  assign new_n1090_ = \a[101]  & \b[101] ;
  assign new_n1091_ = ~new_n1089_ & ~new_n1090_;
  assign new_n1092_ = ~new_n1083_ & ~new_n1087_;
  assign new_n1093_ = ~new_n1091_ & new_n1092_;
  assign new_n1094_ = new_n1091_ & ~new_n1092_;
  assign \f[101]  = ~new_n1093_ & ~new_n1094_;
  assign new_n1096_ = ~\a[102]  & ~\b[102] ;
  assign new_n1097_ = \a[102]  & \b[102] ;
  assign new_n1098_ = ~new_n1096_ & ~new_n1097_;
  assign new_n1099_ = ~new_n1090_ & ~new_n1094_;
  assign new_n1100_ = ~new_n1098_ & new_n1099_;
  assign new_n1101_ = new_n1098_ & ~new_n1099_;
  assign \f[102]  = ~new_n1100_ & ~new_n1101_;
  assign new_n1103_ = ~\a[103]  & ~\b[103] ;
  assign new_n1104_ = \a[103]  & \b[103] ;
  assign new_n1105_ = ~new_n1103_ & ~new_n1104_;
  assign new_n1106_ = ~new_n1097_ & ~new_n1101_;
  assign new_n1107_ = ~new_n1105_ & new_n1106_;
  assign new_n1108_ = new_n1105_ & ~new_n1106_;
  assign \f[103]  = ~new_n1107_ & ~new_n1108_;
  assign new_n1110_ = ~\a[104]  & ~\b[104] ;
  assign new_n1111_ = \a[104]  & \b[104] ;
  assign new_n1112_ = ~new_n1110_ & ~new_n1111_;
  assign new_n1113_ = ~new_n1104_ & ~new_n1108_;
  assign new_n1114_ = ~new_n1112_ & new_n1113_;
  assign new_n1115_ = new_n1112_ & ~new_n1113_;
  assign \f[104]  = ~new_n1114_ & ~new_n1115_;
  assign new_n1117_ = ~\a[105]  & ~\b[105] ;
  assign new_n1118_ = \a[105]  & \b[105] ;
  assign new_n1119_ = ~new_n1117_ & ~new_n1118_;
  assign new_n1120_ = ~new_n1111_ & ~new_n1115_;
  assign new_n1121_ = ~new_n1119_ & new_n1120_;
  assign new_n1122_ = new_n1119_ & ~new_n1120_;
  assign \f[105]  = ~new_n1121_ & ~new_n1122_;
  assign new_n1124_ = ~\a[106]  & ~\b[106] ;
  assign new_n1125_ = \a[106]  & \b[106] ;
  assign new_n1126_ = ~new_n1124_ & ~new_n1125_;
  assign new_n1127_ = ~new_n1118_ & ~new_n1122_;
  assign new_n1128_ = ~new_n1126_ & new_n1127_;
  assign new_n1129_ = new_n1126_ & ~new_n1127_;
  assign \f[106]  = ~new_n1128_ & ~new_n1129_;
  assign new_n1131_ = ~\a[107]  & ~\b[107] ;
  assign new_n1132_ = \a[107]  & \b[107] ;
  assign new_n1133_ = ~new_n1131_ & ~new_n1132_;
  assign new_n1134_ = ~new_n1125_ & ~new_n1129_;
  assign new_n1135_ = ~new_n1133_ & new_n1134_;
  assign new_n1136_ = new_n1133_ & ~new_n1134_;
  assign \f[107]  = ~new_n1135_ & ~new_n1136_;
  assign new_n1138_ = ~\a[108]  & ~\b[108] ;
  assign new_n1139_ = \a[108]  & \b[108] ;
  assign new_n1140_ = ~new_n1138_ & ~new_n1139_;
  assign new_n1141_ = ~new_n1132_ & ~new_n1136_;
  assign new_n1142_ = ~new_n1140_ & new_n1141_;
  assign new_n1143_ = new_n1140_ & ~new_n1141_;
  assign \f[108]  = ~new_n1142_ & ~new_n1143_;
  assign new_n1145_ = ~\a[109]  & ~\b[109] ;
  assign new_n1146_ = \a[109]  & \b[109] ;
  assign new_n1147_ = ~new_n1145_ & ~new_n1146_;
  assign new_n1148_ = ~new_n1139_ & ~new_n1143_;
  assign new_n1149_ = ~new_n1147_ & new_n1148_;
  assign new_n1150_ = new_n1147_ & ~new_n1148_;
  assign \f[109]  = ~new_n1149_ & ~new_n1150_;
  assign new_n1152_ = ~\a[110]  & ~\b[110] ;
  assign new_n1153_ = \a[110]  & \b[110] ;
  assign new_n1154_ = ~new_n1152_ & ~new_n1153_;
  assign new_n1155_ = ~new_n1146_ & ~new_n1150_;
  assign new_n1156_ = ~new_n1154_ & new_n1155_;
  assign new_n1157_ = new_n1154_ & ~new_n1155_;
  assign \f[110]  = ~new_n1156_ & ~new_n1157_;
  assign new_n1159_ = ~\a[111]  & ~\b[111] ;
  assign new_n1160_ = \a[111]  & \b[111] ;
  assign new_n1161_ = ~new_n1159_ & ~new_n1160_;
  assign new_n1162_ = ~new_n1153_ & ~new_n1157_;
  assign new_n1163_ = ~new_n1161_ & new_n1162_;
  assign new_n1164_ = new_n1161_ & ~new_n1162_;
  assign \f[111]  = ~new_n1163_ & ~new_n1164_;
  assign new_n1166_ = ~\a[112]  & ~\b[112] ;
  assign new_n1167_ = \a[112]  & \b[112] ;
  assign new_n1168_ = ~new_n1166_ & ~new_n1167_;
  assign new_n1169_ = ~new_n1160_ & ~new_n1164_;
  assign new_n1170_ = ~new_n1168_ & new_n1169_;
  assign new_n1171_ = new_n1168_ & ~new_n1169_;
  assign \f[112]  = ~new_n1170_ & ~new_n1171_;
  assign new_n1173_ = ~\a[113]  & ~\b[113] ;
  assign new_n1174_ = \a[113]  & \b[113] ;
  assign new_n1175_ = ~new_n1173_ & ~new_n1174_;
  assign new_n1176_ = ~new_n1167_ & ~new_n1171_;
  assign new_n1177_ = ~new_n1175_ & new_n1176_;
  assign new_n1178_ = new_n1175_ & ~new_n1176_;
  assign \f[113]  = ~new_n1177_ & ~new_n1178_;
  assign new_n1180_ = ~\a[114]  & ~\b[114] ;
  assign new_n1181_ = \a[114]  & \b[114] ;
  assign new_n1182_ = ~new_n1180_ & ~new_n1181_;
  assign new_n1183_ = ~new_n1174_ & ~new_n1178_;
  assign new_n1184_ = ~new_n1182_ & new_n1183_;
  assign new_n1185_ = new_n1182_ & ~new_n1183_;
  assign \f[114]  = ~new_n1184_ & ~new_n1185_;
  assign new_n1187_ = ~\a[115]  & ~\b[115] ;
  assign new_n1188_ = \a[115]  & \b[115] ;
  assign new_n1189_ = ~new_n1187_ & ~new_n1188_;
  assign new_n1190_ = ~new_n1181_ & ~new_n1185_;
  assign new_n1191_ = ~new_n1189_ & new_n1190_;
  assign new_n1192_ = new_n1189_ & ~new_n1190_;
  assign \f[115]  = ~new_n1191_ & ~new_n1192_;
  assign new_n1194_ = ~\a[116]  & ~\b[116] ;
  assign new_n1195_ = \a[116]  & \b[116] ;
  assign new_n1196_ = ~new_n1194_ & ~new_n1195_;
  assign new_n1197_ = ~new_n1188_ & ~new_n1192_;
  assign new_n1198_ = ~new_n1196_ & new_n1197_;
  assign new_n1199_ = new_n1196_ & ~new_n1197_;
  assign \f[116]  = ~new_n1198_ & ~new_n1199_;
  assign new_n1201_ = ~\a[117]  & ~\b[117] ;
  assign new_n1202_ = \a[117]  & \b[117] ;
  assign new_n1203_ = ~new_n1201_ & ~new_n1202_;
  assign new_n1204_ = ~new_n1195_ & ~new_n1199_;
  assign new_n1205_ = ~new_n1203_ & new_n1204_;
  assign new_n1206_ = new_n1203_ & ~new_n1204_;
  assign \f[117]  = ~new_n1205_ & ~new_n1206_;
  assign new_n1208_ = ~\a[118]  & ~\b[118] ;
  assign new_n1209_ = \a[118]  & \b[118] ;
  assign new_n1210_ = ~new_n1208_ & ~new_n1209_;
  assign new_n1211_ = ~new_n1202_ & ~new_n1206_;
  assign new_n1212_ = ~new_n1210_ & new_n1211_;
  assign new_n1213_ = new_n1210_ & ~new_n1211_;
  assign \f[118]  = ~new_n1212_ & ~new_n1213_;
  assign new_n1215_ = ~\a[119]  & ~\b[119] ;
  assign new_n1216_ = \a[119]  & \b[119] ;
  assign new_n1217_ = ~new_n1215_ & ~new_n1216_;
  assign new_n1218_ = ~new_n1209_ & ~new_n1213_;
  assign new_n1219_ = ~new_n1217_ & new_n1218_;
  assign new_n1220_ = new_n1217_ & ~new_n1218_;
  assign \f[119]  = ~new_n1219_ & ~new_n1220_;
  assign new_n1222_ = ~\a[120]  & ~\b[120] ;
  assign new_n1223_ = \a[120]  & \b[120] ;
  assign new_n1224_ = ~new_n1222_ & ~new_n1223_;
  assign new_n1225_ = ~new_n1216_ & ~new_n1220_;
  assign new_n1226_ = ~new_n1224_ & new_n1225_;
  assign new_n1227_ = new_n1224_ & ~new_n1225_;
  assign \f[120]  = ~new_n1226_ & ~new_n1227_;
  assign new_n1229_ = ~\a[121]  & ~\b[121] ;
  assign new_n1230_ = \a[121]  & \b[121] ;
  assign new_n1231_ = ~new_n1229_ & ~new_n1230_;
  assign new_n1232_ = ~new_n1223_ & ~new_n1227_;
  assign new_n1233_ = ~new_n1231_ & new_n1232_;
  assign new_n1234_ = new_n1231_ & ~new_n1232_;
  assign \f[121]  = ~new_n1233_ & ~new_n1234_;
  assign new_n1236_ = ~\a[122]  & ~\b[122] ;
  assign new_n1237_ = \a[122]  & \b[122] ;
  assign new_n1238_ = ~new_n1236_ & ~new_n1237_;
  assign new_n1239_ = ~new_n1230_ & ~new_n1234_;
  assign new_n1240_ = ~new_n1238_ & new_n1239_;
  assign new_n1241_ = new_n1238_ & ~new_n1239_;
  assign \f[122]  = ~new_n1240_ & ~new_n1241_;
  assign new_n1243_ = ~\a[123]  & ~\b[123] ;
  assign new_n1244_ = \a[123]  & \b[123] ;
  assign new_n1245_ = ~new_n1243_ & ~new_n1244_;
  assign new_n1246_ = ~new_n1237_ & ~new_n1241_;
  assign new_n1247_ = ~new_n1245_ & new_n1246_;
  assign new_n1248_ = new_n1245_ & ~new_n1246_;
  assign \f[123]  = ~new_n1247_ & ~new_n1248_;
  assign new_n1250_ = ~\a[124]  & ~\b[124] ;
  assign new_n1251_ = \a[124]  & \b[124] ;
  assign new_n1252_ = ~new_n1250_ & ~new_n1251_;
  assign new_n1253_ = ~new_n1244_ & ~new_n1248_;
  assign new_n1254_ = ~new_n1252_ & new_n1253_;
  assign new_n1255_ = new_n1252_ & ~new_n1253_;
  assign \f[124]  = ~new_n1254_ & ~new_n1255_;
  assign new_n1257_ = ~\a[125]  & ~\b[125] ;
  assign new_n1258_ = \a[125]  & \b[125] ;
  assign new_n1259_ = ~new_n1257_ & ~new_n1258_;
  assign new_n1260_ = ~new_n1251_ & ~new_n1255_;
  assign new_n1261_ = ~new_n1259_ & new_n1260_;
  assign new_n1262_ = new_n1259_ & ~new_n1260_;
  assign \f[125]  = ~new_n1261_ & ~new_n1262_;
  assign new_n1264_ = ~\a[126]  & ~\b[126] ;
  assign new_n1265_ = \a[126]  & \b[126] ;
  assign new_n1266_ = ~new_n1264_ & ~new_n1265_;
  assign new_n1267_ = ~new_n1258_ & ~new_n1262_;
  assign new_n1268_ = ~new_n1266_ & new_n1267_;
  assign new_n1269_ = new_n1266_ & ~new_n1267_;
  assign \f[126]  = ~new_n1268_ & ~new_n1269_;
  assign new_n1271_ = ~\a[127]  & ~\b[127] ;
  assign new_n1272_ = \a[127]  & \b[127] ;
  assign new_n1273_ = ~new_n1271_ & ~new_n1272_;
  assign new_n1274_ = ~new_n1265_ & ~new_n1269_;
  assign new_n1275_ = ~new_n1273_ & new_n1274_;
  assign new_n1276_ = new_n1273_ & ~new_n1274_;
  assign \f[127]  = ~new_n1275_ & ~new_n1276_;
  assign cOut = new_n1272_ | new_n1276_;
endmodule



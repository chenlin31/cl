module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128;
  wire n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640;
  assign n257 = x0 & x128;
  assign n258 = (x0 & x128) | (x0 & ~n257) | (x128 & ~n257);
  assign n259 = ~n257 & n258;
  assign n260 = (x1 & x129) | (x1 & n257) | (x129 & n257);
  assign n261 = (~x1 & x129) | (~x1 & n257) | (x129 & n257);
  assign n262 = (x1 & ~n260) | (x1 & n261) | (~n260 & n261);
  assign n263 = (x2 & x130) | (x2 & n260) | (x130 & n260);
  assign n264 = (~x2 & x130) | (~x2 & n260) | (x130 & n260);
  assign n265 = (x2 & ~n263) | (x2 & n264) | (~n263 & n264);
  assign n266 = (x3 & x131) | (x3 & n263) | (x131 & n263);
  assign n267 = (~x3 & x131) | (~x3 & n263) | (x131 & n263);
  assign n268 = (x3 & ~n266) | (x3 & n267) | (~n266 & n267);
  assign n269 = (x4 & x132) | (x4 & n266) | (x132 & n266);
  assign n270 = (~x4 & x132) | (~x4 & n266) | (x132 & n266);
  assign n271 = (x4 & ~n269) | (x4 & n270) | (~n269 & n270);
  assign n272 = (x5 & x133) | (x5 & n269) | (x133 & n269);
  assign n273 = (~x5 & x133) | (~x5 & n269) | (x133 & n269);
  assign n274 = (x5 & ~n272) | (x5 & n273) | (~n272 & n273);
  assign n275 = (x6 & x134) | (x6 & n272) | (x134 & n272);
  assign n276 = (~x6 & x134) | (~x6 & n272) | (x134 & n272);
  assign n277 = (x6 & ~n275) | (x6 & n276) | (~n275 & n276);
  assign n278 = (x7 & x135) | (x7 & n275) | (x135 & n275);
  assign n279 = (~x7 & x135) | (~x7 & n275) | (x135 & n275);
  assign n280 = (x7 & ~n278) | (x7 & n279) | (~n278 & n279);
  assign n281 = (x8 & x136) | (x8 & n278) | (x136 & n278);
  assign n282 = (~x8 & x136) | (~x8 & n278) | (x136 & n278);
  assign n283 = (x8 & ~n281) | (x8 & n282) | (~n281 & n282);
  assign n284 = (x9 & x137) | (x9 & n281) | (x137 & n281);
  assign n285 = (~x9 & x137) | (~x9 & n281) | (x137 & n281);
  assign n286 = (x9 & ~n284) | (x9 & n285) | (~n284 & n285);
  assign n287 = (x10 & x138) | (x10 & n284) | (x138 & n284);
  assign n288 = (~x10 & x138) | (~x10 & n284) | (x138 & n284);
  assign n289 = (x10 & ~n287) | (x10 & n288) | (~n287 & n288);
  assign n290 = (x11 & x139) | (x11 & n287) | (x139 & n287);
  assign n291 = (~x11 & x139) | (~x11 & n287) | (x139 & n287);
  assign n292 = (x11 & ~n290) | (x11 & n291) | (~n290 & n291);
  assign n293 = (x12 & x140) | (x12 & n290) | (x140 & n290);
  assign n294 = (~x12 & x140) | (~x12 & n290) | (x140 & n290);
  assign n295 = (x12 & ~n293) | (x12 & n294) | (~n293 & n294);
  assign n296 = (x13 & x141) | (x13 & n293) | (x141 & n293);
  assign n297 = (~x13 & x141) | (~x13 & n293) | (x141 & n293);
  assign n298 = (x13 & ~n296) | (x13 & n297) | (~n296 & n297);
  assign n299 = (x14 & x142) | (x14 & n296) | (x142 & n296);
  assign n300 = (~x14 & x142) | (~x14 & n296) | (x142 & n296);
  assign n301 = (x14 & ~n299) | (x14 & n300) | (~n299 & n300);
  assign n302 = (x15 & x143) | (x15 & n299) | (x143 & n299);
  assign n303 = (~x15 & x143) | (~x15 & n299) | (x143 & n299);
  assign n304 = (x15 & ~n302) | (x15 & n303) | (~n302 & n303);
  assign n305 = (x16 & x144) | (x16 & n302) | (x144 & n302);
  assign n306 = (~x16 & x144) | (~x16 & n302) | (x144 & n302);
  assign n307 = (x16 & ~n305) | (x16 & n306) | (~n305 & n306);
  assign n308 = (x17 & x145) | (x17 & n305) | (x145 & n305);
  assign n309 = (~x17 & x145) | (~x17 & n305) | (x145 & n305);
  assign n310 = (x17 & ~n308) | (x17 & n309) | (~n308 & n309);
  assign n311 = (x18 & x146) | (x18 & n308) | (x146 & n308);
  assign n312 = (~x18 & x146) | (~x18 & n308) | (x146 & n308);
  assign n313 = (x18 & ~n311) | (x18 & n312) | (~n311 & n312);
  assign n314 = (x19 & x147) | (x19 & n311) | (x147 & n311);
  assign n315 = (~x19 & x147) | (~x19 & n311) | (x147 & n311);
  assign n316 = (x19 & ~n314) | (x19 & n315) | (~n314 & n315);
  assign n317 = (x20 & x148) | (x20 & n314) | (x148 & n314);
  assign n318 = (~x20 & x148) | (~x20 & n314) | (x148 & n314);
  assign n319 = (x20 & ~n317) | (x20 & n318) | (~n317 & n318);
  assign n320 = (x21 & x149) | (x21 & n317) | (x149 & n317);
  assign n321 = (~x21 & x149) | (~x21 & n317) | (x149 & n317);
  assign n322 = (x21 & ~n320) | (x21 & n321) | (~n320 & n321);
  assign n323 = (x22 & x150) | (x22 & n320) | (x150 & n320);
  assign n324 = (~x22 & x150) | (~x22 & n320) | (x150 & n320);
  assign n325 = (x22 & ~n323) | (x22 & n324) | (~n323 & n324);
  assign n326 = (x23 & x151) | (x23 & n323) | (x151 & n323);
  assign n327 = (~x23 & x151) | (~x23 & n323) | (x151 & n323);
  assign n328 = (x23 & ~n326) | (x23 & n327) | (~n326 & n327);
  assign n329 = (x24 & x152) | (x24 & n326) | (x152 & n326);
  assign n330 = (~x24 & x152) | (~x24 & n326) | (x152 & n326);
  assign n331 = (x24 & ~n329) | (x24 & n330) | (~n329 & n330);
  assign n332 = (x25 & x153) | (x25 & n329) | (x153 & n329);
  assign n333 = (~x25 & x153) | (~x25 & n329) | (x153 & n329);
  assign n334 = (x25 & ~n332) | (x25 & n333) | (~n332 & n333);
  assign n335 = (x26 & x154) | (x26 & n332) | (x154 & n332);
  assign n336 = (~x26 & x154) | (~x26 & n332) | (x154 & n332);
  assign n337 = (x26 & ~n335) | (x26 & n336) | (~n335 & n336);
  assign n338 = (x27 & x155) | (x27 & n335) | (x155 & n335);
  assign n339 = (~x27 & x155) | (~x27 & n335) | (x155 & n335);
  assign n340 = (x27 & ~n338) | (x27 & n339) | (~n338 & n339);
  assign n341 = (x28 & x156) | (x28 & n338) | (x156 & n338);
  assign n342 = (~x28 & x156) | (~x28 & n338) | (x156 & n338);
  assign n343 = (x28 & ~n341) | (x28 & n342) | (~n341 & n342);
  assign n344 = (x29 & x157) | (x29 & n341) | (x157 & n341);
  assign n345 = (~x29 & x157) | (~x29 & n341) | (x157 & n341);
  assign n346 = (x29 & ~n344) | (x29 & n345) | (~n344 & n345);
  assign n347 = (x30 & x158) | (x30 & n344) | (x158 & n344);
  assign n348 = (~x30 & x158) | (~x30 & n344) | (x158 & n344);
  assign n349 = (x30 & ~n347) | (x30 & n348) | (~n347 & n348);
  assign n350 = (x31 & x159) | (x31 & n347) | (x159 & n347);
  assign n351 = (~x31 & x159) | (~x31 & n347) | (x159 & n347);
  assign n352 = (x31 & ~n350) | (x31 & n351) | (~n350 & n351);
  assign n353 = (x32 & x160) | (x32 & n350) | (x160 & n350);
  assign n354 = (~x32 & x160) | (~x32 & n350) | (x160 & n350);
  assign n355 = (x32 & ~n353) | (x32 & n354) | (~n353 & n354);
  assign n356 = (x33 & x161) | (x33 & n353) | (x161 & n353);
  assign n357 = (~x33 & x161) | (~x33 & n353) | (x161 & n353);
  assign n358 = (x33 & ~n356) | (x33 & n357) | (~n356 & n357);
  assign n359 = (x34 & x162) | (x34 & n356) | (x162 & n356);
  assign n360 = (~x34 & x162) | (~x34 & n356) | (x162 & n356);
  assign n361 = (x34 & ~n359) | (x34 & n360) | (~n359 & n360);
  assign n362 = (x35 & x163) | (x35 & n359) | (x163 & n359);
  assign n363 = (~x35 & x163) | (~x35 & n359) | (x163 & n359);
  assign n364 = (x35 & ~n362) | (x35 & n363) | (~n362 & n363);
  assign n365 = (x36 & x164) | (x36 & n362) | (x164 & n362);
  assign n366 = (~x36 & x164) | (~x36 & n362) | (x164 & n362);
  assign n367 = (x36 & ~n365) | (x36 & n366) | (~n365 & n366);
  assign n368 = (x37 & x165) | (x37 & n365) | (x165 & n365);
  assign n369 = (~x37 & x165) | (~x37 & n365) | (x165 & n365);
  assign n370 = (x37 & ~n368) | (x37 & n369) | (~n368 & n369);
  assign n371 = (x38 & x166) | (x38 & n368) | (x166 & n368);
  assign n372 = (~x38 & x166) | (~x38 & n368) | (x166 & n368);
  assign n373 = (x38 & ~n371) | (x38 & n372) | (~n371 & n372);
  assign n374 = (x39 & x167) | (x39 & n371) | (x167 & n371);
  assign n375 = (~x39 & x167) | (~x39 & n371) | (x167 & n371);
  assign n376 = (x39 & ~n374) | (x39 & n375) | (~n374 & n375);
  assign n377 = (x40 & x168) | (x40 & n374) | (x168 & n374);
  assign n378 = (~x40 & x168) | (~x40 & n374) | (x168 & n374);
  assign n379 = (x40 & ~n377) | (x40 & n378) | (~n377 & n378);
  assign n380 = (x41 & x169) | (x41 & n377) | (x169 & n377);
  assign n381 = (~x41 & x169) | (~x41 & n377) | (x169 & n377);
  assign n382 = (x41 & ~n380) | (x41 & n381) | (~n380 & n381);
  assign n383 = (x42 & x170) | (x42 & n380) | (x170 & n380);
  assign n384 = (~x42 & x170) | (~x42 & n380) | (x170 & n380);
  assign n385 = (x42 & ~n383) | (x42 & n384) | (~n383 & n384);
  assign n386 = (x43 & x171) | (x43 & n383) | (x171 & n383);
  assign n387 = (~x43 & x171) | (~x43 & n383) | (x171 & n383);
  assign n388 = (x43 & ~n386) | (x43 & n387) | (~n386 & n387);
  assign n389 = (x44 & x172) | (x44 & n386) | (x172 & n386);
  assign n390 = (~x44 & x172) | (~x44 & n386) | (x172 & n386);
  assign n391 = (x44 & ~n389) | (x44 & n390) | (~n389 & n390);
  assign n392 = (x45 & x173) | (x45 & n389) | (x173 & n389);
  assign n393 = (~x45 & x173) | (~x45 & n389) | (x173 & n389);
  assign n394 = (x45 & ~n392) | (x45 & n393) | (~n392 & n393);
  assign n395 = (x46 & x174) | (x46 & n392) | (x174 & n392);
  assign n396 = (~x46 & x174) | (~x46 & n392) | (x174 & n392);
  assign n397 = (x46 & ~n395) | (x46 & n396) | (~n395 & n396);
  assign n398 = (x47 & x175) | (x47 & n395) | (x175 & n395);
  assign n399 = (~x47 & x175) | (~x47 & n395) | (x175 & n395);
  assign n400 = (x47 & ~n398) | (x47 & n399) | (~n398 & n399);
  assign n401 = (x48 & x176) | (x48 & n398) | (x176 & n398);
  assign n402 = (~x48 & x176) | (~x48 & n398) | (x176 & n398);
  assign n403 = (x48 & ~n401) | (x48 & n402) | (~n401 & n402);
  assign n404 = (x49 & x177) | (x49 & n401) | (x177 & n401);
  assign n405 = (~x49 & x177) | (~x49 & n401) | (x177 & n401);
  assign n406 = (x49 & ~n404) | (x49 & n405) | (~n404 & n405);
  assign n407 = (x50 & x178) | (x50 & n404) | (x178 & n404);
  assign n408 = (~x50 & x178) | (~x50 & n404) | (x178 & n404);
  assign n409 = (x50 & ~n407) | (x50 & n408) | (~n407 & n408);
  assign n410 = (x51 & x179) | (x51 & n407) | (x179 & n407);
  assign n411 = (~x51 & x179) | (~x51 & n407) | (x179 & n407);
  assign n412 = (x51 & ~n410) | (x51 & n411) | (~n410 & n411);
  assign n413 = (x52 & x180) | (x52 & n410) | (x180 & n410);
  assign n414 = (~x52 & x180) | (~x52 & n410) | (x180 & n410);
  assign n415 = (x52 & ~n413) | (x52 & n414) | (~n413 & n414);
  assign n416 = (x53 & x181) | (x53 & n413) | (x181 & n413);
  assign n417 = (~x53 & x181) | (~x53 & n413) | (x181 & n413);
  assign n418 = (x53 & ~n416) | (x53 & n417) | (~n416 & n417);
  assign n419 = (x54 & x182) | (x54 & n416) | (x182 & n416);
  assign n420 = (~x54 & x182) | (~x54 & n416) | (x182 & n416);
  assign n421 = (x54 & ~n419) | (x54 & n420) | (~n419 & n420);
  assign n422 = (x55 & x183) | (x55 & n419) | (x183 & n419);
  assign n423 = (~x55 & x183) | (~x55 & n419) | (x183 & n419);
  assign n424 = (x55 & ~n422) | (x55 & n423) | (~n422 & n423);
  assign n425 = (x56 & x184) | (x56 & n422) | (x184 & n422);
  assign n426 = (~x56 & x184) | (~x56 & n422) | (x184 & n422);
  assign n427 = (x56 & ~n425) | (x56 & n426) | (~n425 & n426);
  assign n428 = (x57 & x185) | (x57 & n425) | (x185 & n425);
  assign n429 = (~x57 & x185) | (~x57 & n425) | (x185 & n425);
  assign n430 = (x57 & ~n428) | (x57 & n429) | (~n428 & n429);
  assign n431 = (x58 & x186) | (x58 & n428) | (x186 & n428);
  assign n432 = (~x58 & x186) | (~x58 & n428) | (x186 & n428);
  assign n433 = (x58 & ~n431) | (x58 & n432) | (~n431 & n432);
  assign n434 = (x59 & x187) | (x59 & n431) | (x187 & n431);
  assign n435 = (~x59 & x187) | (~x59 & n431) | (x187 & n431);
  assign n436 = (x59 & ~n434) | (x59 & n435) | (~n434 & n435);
  assign n437 = (x60 & x188) | (x60 & n434) | (x188 & n434);
  assign n438 = (~x60 & x188) | (~x60 & n434) | (x188 & n434);
  assign n439 = (x60 & ~n437) | (x60 & n438) | (~n437 & n438);
  assign n440 = (x61 & x189) | (x61 & n437) | (x189 & n437);
  assign n441 = (~x61 & x189) | (~x61 & n437) | (x189 & n437);
  assign n442 = (x61 & ~n440) | (x61 & n441) | (~n440 & n441);
  assign n443 = (x62 & x190) | (x62 & n440) | (x190 & n440);
  assign n444 = (~x62 & x190) | (~x62 & n440) | (x190 & n440);
  assign n445 = (x62 & ~n443) | (x62 & n444) | (~n443 & n444);
  assign n446 = (x63 & x191) | (x63 & n443) | (x191 & n443);
  assign n447 = (~x63 & x191) | (~x63 & n443) | (x191 & n443);
  assign n448 = (x63 & ~n446) | (x63 & n447) | (~n446 & n447);
  assign n449 = (x64 & x192) | (x64 & n446) | (x192 & n446);
  assign n450 = (~x64 & x192) | (~x64 & n446) | (x192 & n446);
  assign n451 = (x64 & ~n449) | (x64 & n450) | (~n449 & n450);
  assign n452 = (x65 & x193) | (x65 & n449) | (x193 & n449);
  assign n453 = (~x65 & x193) | (~x65 & n449) | (x193 & n449);
  assign n454 = (x65 & ~n452) | (x65 & n453) | (~n452 & n453);
  assign n455 = (x66 & x194) | (x66 & n452) | (x194 & n452);
  assign n456 = (~x66 & x194) | (~x66 & n452) | (x194 & n452);
  assign n457 = (x66 & ~n455) | (x66 & n456) | (~n455 & n456);
  assign n458 = (x67 & x195) | (x67 & n455) | (x195 & n455);
  assign n459 = (~x67 & x195) | (~x67 & n455) | (x195 & n455);
  assign n460 = (x67 & ~n458) | (x67 & n459) | (~n458 & n459);
  assign n461 = (x68 & x196) | (x68 & n458) | (x196 & n458);
  assign n462 = (~x68 & x196) | (~x68 & n458) | (x196 & n458);
  assign n463 = (x68 & ~n461) | (x68 & n462) | (~n461 & n462);
  assign n464 = (x69 & x197) | (x69 & n461) | (x197 & n461);
  assign n465 = (~x69 & x197) | (~x69 & n461) | (x197 & n461);
  assign n466 = (x69 & ~n464) | (x69 & n465) | (~n464 & n465);
  assign n467 = (x70 & x198) | (x70 & n464) | (x198 & n464);
  assign n468 = (~x70 & x198) | (~x70 & n464) | (x198 & n464);
  assign n469 = (x70 & ~n467) | (x70 & n468) | (~n467 & n468);
  assign n470 = (x71 & x199) | (x71 & n467) | (x199 & n467);
  assign n471 = (~x71 & x199) | (~x71 & n467) | (x199 & n467);
  assign n472 = (x71 & ~n470) | (x71 & n471) | (~n470 & n471);
  assign n473 = (x72 & x200) | (x72 & n470) | (x200 & n470);
  assign n474 = (~x72 & x200) | (~x72 & n470) | (x200 & n470);
  assign n475 = (x72 & ~n473) | (x72 & n474) | (~n473 & n474);
  assign n476 = (x73 & x201) | (x73 & n473) | (x201 & n473);
  assign n477 = (~x73 & x201) | (~x73 & n473) | (x201 & n473);
  assign n478 = (x73 & ~n476) | (x73 & n477) | (~n476 & n477);
  assign n479 = (x74 & x202) | (x74 & n476) | (x202 & n476);
  assign n480 = (~x74 & x202) | (~x74 & n476) | (x202 & n476);
  assign n481 = (x74 & ~n479) | (x74 & n480) | (~n479 & n480);
  assign n482 = (x75 & x203) | (x75 & n479) | (x203 & n479);
  assign n483 = (~x75 & x203) | (~x75 & n479) | (x203 & n479);
  assign n484 = (x75 & ~n482) | (x75 & n483) | (~n482 & n483);
  assign n485 = (x76 & x204) | (x76 & n482) | (x204 & n482);
  assign n486 = (~x76 & x204) | (~x76 & n482) | (x204 & n482);
  assign n487 = (x76 & ~n485) | (x76 & n486) | (~n485 & n486);
  assign n488 = (x77 & x205) | (x77 & n485) | (x205 & n485);
  assign n489 = (~x77 & x205) | (~x77 & n485) | (x205 & n485);
  assign n490 = (x77 & ~n488) | (x77 & n489) | (~n488 & n489);
  assign n491 = (x78 & x206) | (x78 & n488) | (x206 & n488);
  assign n492 = (~x78 & x206) | (~x78 & n488) | (x206 & n488);
  assign n493 = (x78 & ~n491) | (x78 & n492) | (~n491 & n492);
  assign n494 = (x79 & x207) | (x79 & n491) | (x207 & n491);
  assign n495 = (~x79 & x207) | (~x79 & n491) | (x207 & n491);
  assign n496 = (x79 & ~n494) | (x79 & n495) | (~n494 & n495);
  assign n497 = (x80 & x208) | (x80 & n494) | (x208 & n494);
  assign n498 = (~x80 & x208) | (~x80 & n494) | (x208 & n494);
  assign n499 = (x80 & ~n497) | (x80 & n498) | (~n497 & n498);
  assign n500 = (x81 & x209) | (x81 & n497) | (x209 & n497);
  assign n501 = (~x81 & x209) | (~x81 & n497) | (x209 & n497);
  assign n502 = (x81 & ~n500) | (x81 & n501) | (~n500 & n501);
  assign n503 = (x82 & x210) | (x82 & n500) | (x210 & n500);
  assign n504 = (~x82 & x210) | (~x82 & n500) | (x210 & n500);
  assign n505 = (x82 & ~n503) | (x82 & n504) | (~n503 & n504);
  assign n506 = (x83 & x211) | (x83 & n503) | (x211 & n503);
  assign n507 = (~x83 & x211) | (~x83 & n503) | (x211 & n503);
  assign n508 = (x83 & ~n506) | (x83 & n507) | (~n506 & n507);
  assign n509 = (x84 & x212) | (x84 & n506) | (x212 & n506);
  assign n510 = (~x84 & x212) | (~x84 & n506) | (x212 & n506);
  assign n511 = (x84 & ~n509) | (x84 & n510) | (~n509 & n510);
  assign n512 = (x85 & x213) | (x85 & n509) | (x213 & n509);
  assign n513 = (~x85 & x213) | (~x85 & n509) | (x213 & n509);
  assign n514 = (x85 & ~n512) | (x85 & n513) | (~n512 & n513);
  assign n515 = (x86 & x214) | (x86 & n512) | (x214 & n512);
  assign n516 = (~x86 & x214) | (~x86 & n512) | (x214 & n512);
  assign n517 = (x86 & ~n515) | (x86 & n516) | (~n515 & n516);
  assign n518 = (x87 & x215) | (x87 & n515) | (x215 & n515);
  assign n519 = (~x87 & x215) | (~x87 & n515) | (x215 & n515);
  assign n520 = (x87 & ~n518) | (x87 & n519) | (~n518 & n519);
  assign n521 = (x88 & x216) | (x88 & n518) | (x216 & n518);
  assign n522 = (~x88 & x216) | (~x88 & n518) | (x216 & n518);
  assign n523 = (x88 & ~n521) | (x88 & n522) | (~n521 & n522);
  assign n524 = (x89 & x217) | (x89 & n521) | (x217 & n521);
  assign n525 = (~x89 & x217) | (~x89 & n521) | (x217 & n521);
  assign n526 = (x89 & ~n524) | (x89 & n525) | (~n524 & n525);
  assign n527 = (x90 & x218) | (x90 & n524) | (x218 & n524);
  assign n528 = (~x90 & x218) | (~x90 & n524) | (x218 & n524);
  assign n529 = (x90 & ~n527) | (x90 & n528) | (~n527 & n528);
  assign n530 = (x91 & x219) | (x91 & n527) | (x219 & n527);
  assign n531 = (~x91 & x219) | (~x91 & n527) | (x219 & n527);
  assign n532 = (x91 & ~n530) | (x91 & n531) | (~n530 & n531);
  assign n533 = (x92 & x220) | (x92 & n530) | (x220 & n530);
  assign n534 = (~x92 & x220) | (~x92 & n530) | (x220 & n530);
  assign n535 = (x92 & ~n533) | (x92 & n534) | (~n533 & n534);
  assign n536 = (x93 & x221) | (x93 & n533) | (x221 & n533);
  assign n537 = (~x93 & x221) | (~x93 & n533) | (x221 & n533);
  assign n538 = (x93 & ~n536) | (x93 & n537) | (~n536 & n537);
  assign n539 = (x94 & x222) | (x94 & n536) | (x222 & n536);
  assign n540 = (~x94 & x222) | (~x94 & n536) | (x222 & n536);
  assign n541 = (x94 & ~n539) | (x94 & n540) | (~n539 & n540);
  assign n542 = (x95 & x223) | (x95 & n539) | (x223 & n539);
  assign n543 = (~x95 & x223) | (~x95 & n539) | (x223 & n539);
  assign n544 = (x95 & ~n542) | (x95 & n543) | (~n542 & n543);
  assign n545 = (x96 & x224) | (x96 & n542) | (x224 & n542);
  assign n546 = (~x96 & x224) | (~x96 & n542) | (x224 & n542);
  assign n547 = (x96 & ~n545) | (x96 & n546) | (~n545 & n546);
  assign n548 = (x97 & x225) | (x97 & n545) | (x225 & n545);
  assign n549 = (~x97 & x225) | (~x97 & n545) | (x225 & n545);
  assign n550 = (x97 & ~n548) | (x97 & n549) | (~n548 & n549);
  assign n551 = (x98 & x226) | (x98 & n548) | (x226 & n548);
  assign n552 = (~x98 & x226) | (~x98 & n548) | (x226 & n548);
  assign n553 = (x98 & ~n551) | (x98 & n552) | (~n551 & n552);
  assign n554 = (x99 & x227) | (x99 & n551) | (x227 & n551);
  assign n555 = (~x99 & x227) | (~x99 & n551) | (x227 & n551);
  assign n556 = (x99 & ~n554) | (x99 & n555) | (~n554 & n555);
  assign n557 = (x100 & x228) | (x100 & n554) | (x228 & n554);
  assign n558 = (~x100 & x228) | (~x100 & n554) | (x228 & n554);
  assign n559 = (x100 & ~n557) | (x100 & n558) | (~n557 & n558);
  assign n560 = (x101 & x229) | (x101 & n557) | (x229 & n557);
  assign n561 = (~x101 & x229) | (~x101 & n557) | (x229 & n557);
  assign n562 = (x101 & ~n560) | (x101 & n561) | (~n560 & n561);
  assign n563 = (x102 & x230) | (x102 & n560) | (x230 & n560);
  assign n564 = (~x102 & x230) | (~x102 & n560) | (x230 & n560);
  assign n565 = (x102 & ~n563) | (x102 & n564) | (~n563 & n564);
  assign n566 = (x103 & x231) | (x103 & n563) | (x231 & n563);
  assign n567 = (~x103 & x231) | (~x103 & n563) | (x231 & n563);
  assign n568 = (x103 & ~n566) | (x103 & n567) | (~n566 & n567);
  assign n569 = (x104 & x232) | (x104 & n566) | (x232 & n566);
  assign n570 = (~x104 & x232) | (~x104 & n566) | (x232 & n566);
  assign n571 = (x104 & ~n569) | (x104 & n570) | (~n569 & n570);
  assign n572 = (x105 & x233) | (x105 & n569) | (x233 & n569);
  assign n573 = (~x105 & x233) | (~x105 & n569) | (x233 & n569);
  assign n574 = (x105 & ~n572) | (x105 & n573) | (~n572 & n573);
  assign n575 = (x106 & x234) | (x106 & n572) | (x234 & n572);
  assign n576 = (~x106 & x234) | (~x106 & n572) | (x234 & n572);
  assign n577 = (x106 & ~n575) | (x106 & n576) | (~n575 & n576);
  assign n578 = (x107 & x235) | (x107 & n575) | (x235 & n575);
  assign n579 = (~x107 & x235) | (~x107 & n575) | (x235 & n575);
  assign n580 = (x107 & ~n578) | (x107 & n579) | (~n578 & n579);
  assign n581 = (x108 & x236) | (x108 & n578) | (x236 & n578);
  assign n582 = (~x108 & x236) | (~x108 & n578) | (x236 & n578);
  assign n583 = (x108 & ~n581) | (x108 & n582) | (~n581 & n582);
  assign n584 = (x109 & x237) | (x109 & n581) | (x237 & n581);
  assign n585 = (~x109 & x237) | (~x109 & n581) | (x237 & n581);
  assign n586 = (x109 & ~n584) | (x109 & n585) | (~n584 & n585);
  assign n587 = (x110 & x238) | (x110 & n584) | (x238 & n584);
  assign n588 = (~x110 & x238) | (~x110 & n584) | (x238 & n584);
  assign n589 = (x110 & ~n587) | (x110 & n588) | (~n587 & n588);
  assign n590 = (x111 & x239) | (x111 & n587) | (x239 & n587);
  assign n591 = (~x111 & x239) | (~x111 & n587) | (x239 & n587);
  assign n592 = (x111 & ~n590) | (x111 & n591) | (~n590 & n591);
  assign n593 = (x112 & x240) | (x112 & n590) | (x240 & n590);
  assign n594 = (~x112 & x240) | (~x112 & n590) | (x240 & n590);
  assign n595 = (x112 & ~n593) | (x112 & n594) | (~n593 & n594);
  assign n596 = (x113 & x241) | (x113 & n593) | (x241 & n593);
  assign n597 = (~x113 & x241) | (~x113 & n593) | (x241 & n593);
  assign n598 = (x113 & ~n596) | (x113 & n597) | (~n596 & n597);
  assign n599 = (x114 & x242) | (x114 & n596) | (x242 & n596);
  assign n600 = (~x114 & x242) | (~x114 & n596) | (x242 & n596);
  assign n601 = (x114 & ~n599) | (x114 & n600) | (~n599 & n600);
  assign n602 = (x115 & x243) | (x115 & n599) | (x243 & n599);
  assign n603 = (~x115 & x243) | (~x115 & n599) | (x243 & n599);
  assign n604 = (x115 & ~n602) | (x115 & n603) | (~n602 & n603);
  assign n605 = (x116 & x244) | (x116 & n602) | (x244 & n602);
  assign n606 = (~x116 & x244) | (~x116 & n602) | (x244 & n602);
  assign n607 = (x116 & ~n605) | (x116 & n606) | (~n605 & n606);
  assign n608 = (x117 & x245) | (x117 & n605) | (x245 & n605);
  assign n609 = (~x117 & x245) | (~x117 & n605) | (x245 & n605);
  assign n610 = (x117 & ~n608) | (x117 & n609) | (~n608 & n609);
  assign n611 = (x118 & x246) | (x118 & n608) | (x246 & n608);
  assign n612 = (~x118 & x246) | (~x118 & n608) | (x246 & n608);
  assign n613 = (x118 & ~n611) | (x118 & n612) | (~n611 & n612);
  assign n614 = (x119 & x247) | (x119 & n611) | (x247 & n611);
  assign n615 = (~x119 & x247) | (~x119 & n611) | (x247 & n611);
  assign n616 = (x119 & ~n614) | (x119 & n615) | (~n614 & n615);
  assign n617 = (x120 & x248) | (x120 & n614) | (x248 & n614);
  assign n618 = (~x120 & x248) | (~x120 & n614) | (x248 & n614);
  assign n619 = (x120 & ~n617) | (x120 & n618) | (~n617 & n618);
  assign n620 = (x121 & x249) | (x121 & n617) | (x249 & n617);
  assign n621 = (~x121 & x249) | (~x121 & n617) | (x249 & n617);
  assign n622 = (x121 & ~n620) | (x121 & n621) | (~n620 & n621);
  assign n623 = (x122 & x250) | (x122 & n620) | (x250 & n620);
  assign n624 = (~x122 & x250) | (~x122 & n620) | (x250 & n620);
  assign n625 = (x122 & ~n623) | (x122 & n624) | (~n623 & n624);
  assign n626 = (x123 & x251) | (x123 & n623) | (x251 & n623);
  assign n627 = (~x123 & x251) | (~x123 & n623) | (x251 & n623);
  assign n628 = (x123 & ~n626) | (x123 & n627) | (~n626 & n627);
  assign n629 = (x124 & x252) | (x124 & n626) | (x252 & n626);
  assign n630 = (~x124 & x252) | (~x124 & n626) | (x252 & n626);
  assign n631 = (x124 & ~n629) | (x124 & n630) | (~n629 & n630);
  assign n632 = (x125 & x253) | (x125 & n629) | (x253 & n629);
  assign n633 = (~x125 & x253) | (~x125 & n629) | (x253 & n629);
  assign n634 = (x125 & ~n632) | (x125 & n633) | (~n632 & n633);
  assign n635 = (x126 & x254) | (x126 & n632) | (x254 & n632);
  assign n636 = (~x126 & x254) | (~x126 & n632) | (x254 & n632);
  assign n637 = (x126 & ~n635) | (x126 & n636) | (~n635 & n636);
  assign n638 = (x127 & x255) | (x127 & n635) | (x255 & n635);
  assign n639 = (~x127 & x255) | (~x127 & n635) | (x255 & n635);
  assign n640 = (x127 & ~n638) | (x127 & n639) | (~n638 & n639);
  assign y0 = n259;
  assign y1 = n262;
  assign y2 = n265;
  assign y3 = n268;
  assign y4 = n271;
  assign y5 = n274;
  assign y6 = n277;
  assign y7 = n280;
  assign y8 = n283;
  assign y9 = n286;
  assign y10 = n289;
  assign y11 = n292;
  assign y12 = n295;
  assign y13 = n298;
  assign y14 = n301;
  assign y15 = n304;
  assign y16 = n307;
  assign y17 = n310;
  assign y18 = n313;
  assign y19 = n316;
  assign y20 = n319;
  assign y21 = n322;
  assign y22 = n325;
  assign y23 = n328;
  assign y24 = n331;
  assign y25 = n334;
  assign y26 = n337;
  assign y27 = n340;
  assign y28 = n343;
  assign y29 = n346;
  assign y30 = n349;
  assign y31 = n352;
  assign y32 = n355;
  assign y33 = n358;
  assign y34 = n361;
  assign y35 = n364;
  assign y36 = n367;
  assign y37 = n370;
  assign y38 = n373;
  assign y39 = n376;
  assign y40 = n379;
  assign y41 = n382;
  assign y42 = n385;
  assign y43 = n388;
  assign y44 = n391;
  assign y45 = n394;
  assign y46 = n397;
  assign y47 = n400;
  assign y48 = n403;
  assign y49 = n406;
  assign y50 = n409;
  assign y51 = n412;
  assign y52 = n415;
  assign y53 = n418;
  assign y54 = n421;
  assign y55 = n424;
  assign y56 = n427;
  assign y57 = n430;
  assign y58 = n433;
  assign y59 = n436;
  assign y60 = n439;
  assign y61 = n442;
  assign y62 = n445;
  assign y63 = n448;
  assign y64 = n451;
  assign y65 = n454;
  assign y66 = n457;
  assign y67 = n460;
  assign y68 = n463;
  assign y69 = n466;
  assign y70 = n469;
  assign y71 = n472;
  assign y72 = n475;
  assign y73 = n478;
  assign y74 = n481;
  assign y75 = n484;
  assign y76 = n487;
  assign y77 = n490;
  assign y78 = n493;
  assign y79 = n496;
  assign y80 = n499;
  assign y81 = n502;
  assign y82 = n505;
  assign y83 = n508;
  assign y84 = n511;
  assign y85 = n514;
  assign y86 = n517;
  assign y87 = n520;
  assign y88 = n523;
  assign y89 = n526;
  assign y90 = n529;
  assign y91 = n532;
  assign y92 = n535;
  assign y93 = n538;
  assign y94 = n541;
  assign y95 = n544;
  assign y96 = n547;
  assign y97 = n550;
  assign y98 = n553;
  assign y99 = n556;
  assign y100 = n559;
  assign y101 = n562;
  assign y102 = n565;
  assign y103 = n568;
  assign y104 = n571;
  assign y105 = n574;
  assign y106 = n577;
  assign y107 = n580;
  assign y108 = n583;
  assign y109 = n586;
  assign y110 = n589;
  assign y111 = n592;
  assign y112 = n595;
  assign y113 = n598;
  assign y114 = n601;
  assign y115 = n604;
  assign y116 = n607;
  assign y117 = n610;
  assign y118 = n613;
  assign y119 = n616;
  assign y120 = n619;
  assign y121 = n622;
  assign y122 = n625;
  assign y123 = n628;
  assign y124 = n631;
  assign y125 = n634;
  assign y126 = n637;
  assign y127 = n640;
  assign y128 = n638;
endmodule
